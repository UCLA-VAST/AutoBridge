module kernel0_kernel0_ap_fadd_5_full_dsp_32 (
    input aclk                 ,
    input aclken               ,
    input s_axis_a_tvalid      ,
    input s_axis_a_tdata       ,
    input s_axis_b_tvalid      ,
    input s_axis_b_tdata       ,
    output m_axis_result_tvalid ,
    output m_axis_result_tdata  
);

endmodule