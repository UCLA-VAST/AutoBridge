`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO = "PageRank_PageRank,hls_ip_2019_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcu280-fsvh2892-2L-e,HLS_INPUT_CLOCK=4.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=1,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=1460,HLS_SYN_LUT=2647,HLS_VERSION=2019_2}" *)


module PageRank
(
  ap_clk,
  ap_rst_n,
  s_axi_control_AWVALID,
  s_axi_control_AWREADY,
  s_axi_control_AWADDR,
  s_axi_control_WVALID,
  s_axi_control_WREADY,
  s_axi_control_WDATA,
  s_axi_control_WSTRB,
  s_axi_control_ARVALID,
  s_axi_control_ARREADY,
  s_axi_control_ARADDR,
  s_axi_control_RVALID,
  s_axi_control_RREADY,
  s_axi_control_RDATA,
  s_axi_control_RRESP,
  s_axi_control_BVALID,
  s_axi_control_BREADY,
  s_axi_control_BRESP,
  interrupt,
  m_axi_metadata_ARADDR,
  m_axi_metadata_ARBURST,
  m_axi_metadata_ARCACHE,
  m_axi_metadata_ARID,
  m_axi_metadata_ARLEN,
  m_axi_metadata_ARLOCK,
  m_axi_metadata_ARPROT,
  m_axi_metadata_ARQOS,
  m_axi_metadata_ARREADY,
  m_axi_metadata_ARREGION,
  m_axi_metadata_ARSIZE,
  m_axi_metadata_ARUSER,
  m_axi_metadata_ARVALID,
  m_axi_metadata_AWADDR,
  m_axi_metadata_AWBURST,
  m_axi_metadata_AWCACHE,
  m_axi_metadata_AWID,
  m_axi_metadata_AWLEN,
  m_axi_metadata_AWLOCK,
  m_axi_metadata_AWPROT,
  m_axi_metadata_AWQOS,
  m_axi_metadata_AWREADY,
  m_axi_metadata_AWREGION,
  m_axi_metadata_AWSIZE,
  m_axi_metadata_AWUSER,
  m_axi_metadata_AWVALID,
  m_axi_metadata_BID,
  m_axi_metadata_BREADY,
  m_axi_metadata_BRESP,
  m_axi_metadata_BUSER,
  m_axi_metadata_BVALID,
  m_axi_metadata_RDATA,
  m_axi_metadata_RID,
  m_axi_metadata_RLAST,
  m_axi_metadata_RREADY,
  m_axi_metadata_RRESP,
  m_axi_metadata_RUSER,
  m_axi_metadata_RVALID,
  m_axi_metadata_WDATA,
  m_axi_metadata_WID,
  m_axi_metadata_WLAST,
  m_axi_metadata_WREADY,
  m_axi_metadata_WSTRB,
  m_axi_metadata_WUSER,
  m_axi_metadata_WVALID,
  m_axi_edges_0_ARADDR,
  m_axi_edges_0_ARBURST,
  m_axi_edges_0_ARCACHE,
  m_axi_edges_0_ARID,
  m_axi_edges_0_ARLEN,
  m_axi_edges_0_ARLOCK,
  m_axi_edges_0_ARPROT,
  m_axi_edges_0_ARQOS,
  m_axi_edges_0_ARREADY,
  m_axi_edges_0_ARREGION,
  m_axi_edges_0_ARSIZE,
  m_axi_edges_0_ARUSER,
  m_axi_edges_0_ARVALID,
  m_axi_edges_0_AWADDR,
  m_axi_edges_0_AWBURST,
  m_axi_edges_0_AWCACHE,
  m_axi_edges_0_AWID,
  m_axi_edges_0_AWLEN,
  m_axi_edges_0_AWLOCK,
  m_axi_edges_0_AWPROT,
  m_axi_edges_0_AWQOS,
  m_axi_edges_0_AWREADY,
  m_axi_edges_0_AWREGION,
  m_axi_edges_0_AWSIZE,
  m_axi_edges_0_AWUSER,
  m_axi_edges_0_AWVALID,
  m_axi_edges_0_BID,
  m_axi_edges_0_BREADY,
  m_axi_edges_0_BRESP,
  m_axi_edges_0_BUSER,
  m_axi_edges_0_BVALID,
  m_axi_edges_0_RDATA,
  m_axi_edges_0_RID,
  m_axi_edges_0_RLAST,
  m_axi_edges_0_RREADY,
  m_axi_edges_0_RRESP,
  m_axi_edges_0_RUSER,
  m_axi_edges_0_RVALID,
  m_axi_edges_0_WDATA,
  m_axi_edges_0_WID,
  m_axi_edges_0_WLAST,
  m_axi_edges_0_WREADY,
  m_axi_edges_0_WSTRB,
  m_axi_edges_0_WUSER,
  m_axi_edges_0_WVALID,
  m_axi_edges_1_ARADDR,
  m_axi_edges_1_ARBURST,
  m_axi_edges_1_ARCACHE,
  m_axi_edges_1_ARID,
  m_axi_edges_1_ARLEN,
  m_axi_edges_1_ARLOCK,
  m_axi_edges_1_ARPROT,
  m_axi_edges_1_ARQOS,
  m_axi_edges_1_ARREADY,
  m_axi_edges_1_ARREGION,
  m_axi_edges_1_ARSIZE,
  m_axi_edges_1_ARUSER,
  m_axi_edges_1_ARVALID,
  m_axi_edges_1_AWADDR,
  m_axi_edges_1_AWBURST,
  m_axi_edges_1_AWCACHE,
  m_axi_edges_1_AWID,
  m_axi_edges_1_AWLEN,
  m_axi_edges_1_AWLOCK,
  m_axi_edges_1_AWPROT,
  m_axi_edges_1_AWQOS,
  m_axi_edges_1_AWREADY,
  m_axi_edges_1_AWREGION,
  m_axi_edges_1_AWSIZE,
  m_axi_edges_1_AWUSER,
  m_axi_edges_1_AWVALID,
  m_axi_edges_1_BID,
  m_axi_edges_1_BREADY,
  m_axi_edges_1_BRESP,
  m_axi_edges_1_BUSER,
  m_axi_edges_1_BVALID,
  m_axi_edges_1_RDATA,
  m_axi_edges_1_RID,
  m_axi_edges_1_RLAST,
  m_axi_edges_1_RREADY,
  m_axi_edges_1_RRESP,
  m_axi_edges_1_RUSER,
  m_axi_edges_1_RVALID,
  m_axi_edges_1_WDATA,
  m_axi_edges_1_WID,
  m_axi_edges_1_WLAST,
  m_axi_edges_1_WREADY,
  m_axi_edges_1_WSTRB,
  m_axi_edges_1_WUSER,
  m_axi_edges_1_WVALID,
  m_axi_edges_2_ARADDR,
  m_axi_edges_2_ARBURST,
  m_axi_edges_2_ARCACHE,
  m_axi_edges_2_ARID,
  m_axi_edges_2_ARLEN,
  m_axi_edges_2_ARLOCK,
  m_axi_edges_2_ARPROT,
  m_axi_edges_2_ARQOS,
  m_axi_edges_2_ARREADY,
  m_axi_edges_2_ARREGION,
  m_axi_edges_2_ARSIZE,
  m_axi_edges_2_ARUSER,
  m_axi_edges_2_ARVALID,
  m_axi_edges_2_AWADDR,
  m_axi_edges_2_AWBURST,
  m_axi_edges_2_AWCACHE,
  m_axi_edges_2_AWID,
  m_axi_edges_2_AWLEN,
  m_axi_edges_2_AWLOCK,
  m_axi_edges_2_AWPROT,
  m_axi_edges_2_AWQOS,
  m_axi_edges_2_AWREADY,
  m_axi_edges_2_AWREGION,
  m_axi_edges_2_AWSIZE,
  m_axi_edges_2_AWUSER,
  m_axi_edges_2_AWVALID,
  m_axi_edges_2_BID,
  m_axi_edges_2_BREADY,
  m_axi_edges_2_BRESP,
  m_axi_edges_2_BUSER,
  m_axi_edges_2_BVALID,
  m_axi_edges_2_RDATA,
  m_axi_edges_2_RID,
  m_axi_edges_2_RLAST,
  m_axi_edges_2_RREADY,
  m_axi_edges_2_RRESP,
  m_axi_edges_2_RUSER,
  m_axi_edges_2_RVALID,
  m_axi_edges_2_WDATA,
  m_axi_edges_2_WID,
  m_axi_edges_2_WLAST,
  m_axi_edges_2_WREADY,
  m_axi_edges_2_WSTRB,
  m_axi_edges_2_WUSER,
  m_axi_edges_2_WVALID,
  m_axi_edges_3_ARADDR,
  m_axi_edges_3_ARBURST,
  m_axi_edges_3_ARCACHE,
  m_axi_edges_3_ARID,
  m_axi_edges_3_ARLEN,
  m_axi_edges_3_ARLOCK,
  m_axi_edges_3_ARPROT,
  m_axi_edges_3_ARQOS,
  m_axi_edges_3_ARREADY,
  m_axi_edges_3_ARREGION,
  m_axi_edges_3_ARSIZE,
  m_axi_edges_3_ARUSER,
  m_axi_edges_3_ARVALID,
  m_axi_edges_3_AWADDR,
  m_axi_edges_3_AWBURST,
  m_axi_edges_3_AWCACHE,
  m_axi_edges_3_AWID,
  m_axi_edges_3_AWLEN,
  m_axi_edges_3_AWLOCK,
  m_axi_edges_3_AWPROT,
  m_axi_edges_3_AWQOS,
  m_axi_edges_3_AWREADY,
  m_axi_edges_3_AWREGION,
  m_axi_edges_3_AWSIZE,
  m_axi_edges_3_AWUSER,
  m_axi_edges_3_AWVALID,
  m_axi_edges_3_BID,
  m_axi_edges_3_BREADY,
  m_axi_edges_3_BRESP,
  m_axi_edges_3_BUSER,
  m_axi_edges_3_BVALID,
  m_axi_edges_3_RDATA,
  m_axi_edges_3_RID,
  m_axi_edges_3_RLAST,
  m_axi_edges_3_RREADY,
  m_axi_edges_3_RRESP,
  m_axi_edges_3_RUSER,
  m_axi_edges_3_RVALID,
  m_axi_edges_3_WDATA,
  m_axi_edges_3_WID,
  m_axi_edges_3_WLAST,
  m_axi_edges_3_WREADY,
  m_axi_edges_3_WSTRB,
  m_axi_edges_3_WUSER,
  m_axi_edges_3_WVALID,
  m_axi_edges_4_ARADDR,
  m_axi_edges_4_ARBURST,
  m_axi_edges_4_ARCACHE,
  m_axi_edges_4_ARID,
  m_axi_edges_4_ARLEN,
  m_axi_edges_4_ARLOCK,
  m_axi_edges_4_ARPROT,
  m_axi_edges_4_ARQOS,
  m_axi_edges_4_ARREADY,
  m_axi_edges_4_ARREGION,
  m_axi_edges_4_ARSIZE,
  m_axi_edges_4_ARUSER,
  m_axi_edges_4_ARVALID,
  m_axi_edges_4_AWADDR,
  m_axi_edges_4_AWBURST,
  m_axi_edges_4_AWCACHE,
  m_axi_edges_4_AWID,
  m_axi_edges_4_AWLEN,
  m_axi_edges_4_AWLOCK,
  m_axi_edges_4_AWPROT,
  m_axi_edges_4_AWQOS,
  m_axi_edges_4_AWREADY,
  m_axi_edges_4_AWREGION,
  m_axi_edges_4_AWSIZE,
  m_axi_edges_4_AWUSER,
  m_axi_edges_4_AWVALID,
  m_axi_edges_4_BID,
  m_axi_edges_4_BREADY,
  m_axi_edges_4_BRESP,
  m_axi_edges_4_BUSER,
  m_axi_edges_4_BVALID,
  m_axi_edges_4_RDATA,
  m_axi_edges_4_RID,
  m_axi_edges_4_RLAST,
  m_axi_edges_4_RREADY,
  m_axi_edges_4_RRESP,
  m_axi_edges_4_RUSER,
  m_axi_edges_4_RVALID,
  m_axi_edges_4_WDATA,
  m_axi_edges_4_WID,
  m_axi_edges_4_WLAST,
  m_axi_edges_4_WREADY,
  m_axi_edges_4_WSTRB,
  m_axi_edges_4_WUSER,
  m_axi_edges_4_WVALID,
  m_axi_edges_5_ARADDR,
  m_axi_edges_5_ARBURST,
  m_axi_edges_5_ARCACHE,
  m_axi_edges_5_ARID,
  m_axi_edges_5_ARLEN,
  m_axi_edges_5_ARLOCK,
  m_axi_edges_5_ARPROT,
  m_axi_edges_5_ARQOS,
  m_axi_edges_5_ARREADY,
  m_axi_edges_5_ARREGION,
  m_axi_edges_5_ARSIZE,
  m_axi_edges_5_ARUSER,
  m_axi_edges_5_ARVALID,
  m_axi_edges_5_AWADDR,
  m_axi_edges_5_AWBURST,
  m_axi_edges_5_AWCACHE,
  m_axi_edges_5_AWID,
  m_axi_edges_5_AWLEN,
  m_axi_edges_5_AWLOCK,
  m_axi_edges_5_AWPROT,
  m_axi_edges_5_AWQOS,
  m_axi_edges_5_AWREADY,
  m_axi_edges_5_AWREGION,
  m_axi_edges_5_AWSIZE,
  m_axi_edges_5_AWUSER,
  m_axi_edges_5_AWVALID,
  m_axi_edges_5_BID,
  m_axi_edges_5_BREADY,
  m_axi_edges_5_BRESP,
  m_axi_edges_5_BUSER,
  m_axi_edges_5_BVALID,
  m_axi_edges_5_RDATA,
  m_axi_edges_5_RID,
  m_axi_edges_5_RLAST,
  m_axi_edges_5_RREADY,
  m_axi_edges_5_RRESP,
  m_axi_edges_5_RUSER,
  m_axi_edges_5_RVALID,
  m_axi_edges_5_WDATA,
  m_axi_edges_5_WID,
  m_axi_edges_5_WLAST,
  m_axi_edges_5_WREADY,
  m_axi_edges_5_WSTRB,
  m_axi_edges_5_WUSER,
  m_axi_edges_5_WVALID,
  m_axi_edges_6_ARADDR,
  m_axi_edges_6_ARBURST,
  m_axi_edges_6_ARCACHE,
  m_axi_edges_6_ARID,
  m_axi_edges_6_ARLEN,
  m_axi_edges_6_ARLOCK,
  m_axi_edges_6_ARPROT,
  m_axi_edges_6_ARQOS,
  m_axi_edges_6_ARREADY,
  m_axi_edges_6_ARREGION,
  m_axi_edges_6_ARSIZE,
  m_axi_edges_6_ARUSER,
  m_axi_edges_6_ARVALID,
  m_axi_edges_6_AWADDR,
  m_axi_edges_6_AWBURST,
  m_axi_edges_6_AWCACHE,
  m_axi_edges_6_AWID,
  m_axi_edges_6_AWLEN,
  m_axi_edges_6_AWLOCK,
  m_axi_edges_6_AWPROT,
  m_axi_edges_6_AWQOS,
  m_axi_edges_6_AWREADY,
  m_axi_edges_6_AWREGION,
  m_axi_edges_6_AWSIZE,
  m_axi_edges_6_AWUSER,
  m_axi_edges_6_AWVALID,
  m_axi_edges_6_BID,
  m_axi_edges_6_BREADY,
  m_axi_edges_6_BRESP,
  m_axi_edges_6_BUSER,
  m_axi_edges_6_BVALID,
  m_axi_edges_6_RDATA,
  m_axi_edges_6_RID,
  m_axi_edges_6_RLAST,
  m_axi_edges_6_RREADY,
  m_axi_edges_6_RRESP,
  m_axi_edges_6_RUSER,
  m_axi_edges_6_RVALID,
  m_axi_edges_6_WDATA,
  m_axi_edges_6_WID,
  m_axi_edges_6_WLAST,
  m_axi_edges_6_WREADY,
  m_axi_edges_6_WSTRB,
  m_axi_edges_6_WUSER,
  m_axi_edges_6_WVALID,
  m_axi_edges_7_ARADDR,
  m_axi_edges_7_ARBURST,
  m_axi_edges_7_ARCACHE,
  m_axi_edges_7_ARID,
  m_axi_edges_7_ARLEN,
  m_axi_edges_7_ARLOCK,
  m_axi_edges_7_ARPROT,
  m_axi_edges_7_ARQOS,
  m_axi_edges_7_ARREADY,
  m_axi_edges_7_ARREGION,
  m_axi_edges_7_ARSIZE,
  m_axi_edges_7_ARUSER,
  m_axi_edges_7_ARVALID,
  m_axi_edges_7_AWADDR,
  m_axi_edges_7_AWBURST,
  m_axi_edges_7_AWCACHE,
  m_axi_edges_7_AWID,
  m_axi_edges_7_AWLEN,
  m_axi_edges_7_AWLOCK,
  m_axi_edges_7_AWPROT,
  m_axi_edges_7_AWQOS,
  m_axi_edges_7_AWREADY,
  m_axi_edges_7_AWREGION,
  m_axi_edges_7_AWSIZE,
  m_axi_edges_7_AWUSER,
  m_axi_edges_7_AWVALID,
  m_axi_edges_7_BID,
  m_axi_edges_7_BREADY,
  m_axi_edges_7_BRESP,
  m_axi_edges_7_BUSER,
  m_axi_edges_7_BVALID,
  m_axi_edges_7_RDATA,
  m_axi_edges_7_RID,
  m_axi_edges_7_RLAST,
  m_axi_edges_7_RREADY,
  m_axi_edges_7_RRESP,
  m_axi_edges_7_RUSER,
  m_axi_edges_7_RVALID,
  m_axi_edges_7_WDATA,
  m_axi_edges_7_WID,
  m_axi_edges_7_WLAST,
  m_axi_edges_7_WREADY,
  m_axi_edges_7_WSTRB,
  m_axi_edges_7_WUSER,
  m_axi_edges_7_WVALID,
  m_axi_updates_0_ARADDR,
  m_axi_updates_0_ARBURST,
  m_axi_updates_0_ARCACHE,
  m_axi_updates_0_ARID,
  m_axi_updates_0_ARLEN,
  m_axi_updates_0_ARLOCK,
  m_axi_updates_0_ARPROT,
  m_axi_updates_0_ARQOS,
  m_axi_updates_0_ARREADY,
  m_axi_updates_0_ARREGION,
  m_axi_updates_0_ARSIZE,
  m_axi_updates_0_ARUSER,
  m_axi_updates_0_ARVALID,
  m_axi_updates_0_AWADDR,
  m_axi_updates_0_AWBURST,
  m_axi_updates_0_AWCACHE,
  m_axi_updates_0_AWID,
  m_axi_updates_0_AWLEN,
  m_axi_updates_0_AWLOCK,
  m_axi_updates_0_AWPROT,
  m_axi_updates_0_AWQOS,
  m_axi_updates_0_AWREADY,
  m_axi_updates_0_AWREGION,
  m_axi_updates_0_AWSIZE,
  m_axi_updates_0_AWUSER,
  m_axi_updates_0_AWVALID,
  m_axi_updates_0_BID,
  m_axi_updates_0_BREADY,
  m_axi_updates_0_BRESP,
  m_axi_updates_0_BUSER,
  m_axi_updates_0_BVALID,
  m_axi_updates_0_RDATA,
  m_axi_updates_0_RID,
  m_axi_updates_0_RLAST,
  m_axi_updates_0_RREADY,
  m_axi_updates_0_RRESP,
  m_axi_updates_0_RUSER,
  m_axi_updates_0_RVALID,
  m_axi_updates_0_WDATA,
  m_axi_updates_0_WID,
  m_axi_updates_0_WLAST,
  m_axi_updates_0_WREADY,
  m_axi_updates_0_WSTRB,
  m_axi_updates_0_WUSER,
  m_axi_updates_0_WVALID,
  m_axi_updates_1_ARADDR,
  m_axi_updates_1_ARBURST,
  m_axi_updates_1_ARCACHE,
  m_axi_updates_1_ARID,
  m_axi_updates_1_ARLEN,
  m_axi_updates_1_ARLOCK,
  m_axi_updates_1_ARPROT,
  m_axi_updates_1_ARQOS,
  m_axi_updates_1_ARREADY,
  m_axi_updates_1_ARREGION,
  m_axi_updates_1_ARSIZE,
  m_axi_updates_1_ARUSER,
  m_axi_updates_1_ARVALID,
  m_axi_updates_1_AWADDR,
  m_axi_updates_1_AWBURST,
  m_axi_updates_1_AWCACHE,
  m_axi_updates_1_AWID,
  m_axi_updates_1_AWLEN,
  m_axi_updates_1_AWLOCK,
  m_axi_updates_1_AWPROT,
  m_axi_updates_1_AWQOS,
  m_axi_updates_1_AWREADY,
  m_axi_updates_1_AWREGION,
  m_axi_updates_1_AWSIZE,
  m_axi_updates_1_AWUSER,
  m_axi_updates_1_AWVALID,
  m_axi_updates_1_BID,
  m_axi_updates_1_BREADY,
  m_axi_updates_1_BRESP,
  m_axi_updates_1_BUSER,
  m_axi_updates_1_BVALID,
  m_axi_updates_1_RDATA,
  m_axi_updates_1_RID,
  m_axi_updates_1_RLAST,
  m_axi_updates_1_RREADY,
  m_axi_updates_1_RRESP,
  m_axi_updates_1_RUSER,
  m_axi_updates_1_RVALID,
  m_axi_updates_1_WDATA,
  m_axi_updates_1_WID,
  m_axi_updates_1_WLAST,
  m_axi_updates_1_WREADY,
  m_axi_updates_1_WSTRB,
  m_axi_updates_1_WUSER,
  m_axi_updates_1_WVALID,
  m_axi_updates_2_ARADDR,
  m_axi_updates_2_ARBURST,
  m_axi_updates_2_ARCACHE,
  m_axi_updates_2_ARID,
  m_axi_updates_2_ARLEN,
  m_axi_updates_2_ARLOCK,
  m_axi_updates_2_ARPROT,
  m_axi_updates_2_ARQOS,
  m_axi_updates_2_ARREADY,
  m_axi_updates_2_ARREGION,
  m_axi_updates_2_ARSIZE,
  m_axi_updates_2_ARUSER,
  m_axi_updates_2_ARVALID,
  m_axi_updates_2_AWADDR,
  m_axi_updates_2_AWBURST,
  m_axi_updates_2_AWCACHE,
  m_axi_updates_2_AWID,
  m_axi_updates_2_AWLEN,
  m_axi_updates_2_AWLOCK,
  m_axi_updates_2_AWPROT,
  m_axi_updates_2_AWQOS,
  m_axi_updates_2_AWREADY,
  m_axi_updates_2_AWREGION,
  m_axi_updates_2_AWSIZE,
  m_axi_updates_2_AWUSER,
  m_axi_updates_2_AWVALID,
  m_axi_updates_2_BID,
  m_axi_updates_2_BREADY,
  m_axi_updates_2_BRESP,
  m_axi_updates_2_BUSER,
  m_axi_updates_2_BVALID,
  m_axi_updates_2_RDATA,
  m_axi_updates_2_RID,
  m_axi_updates_2_RLAST,
  m_axi_updates_2_RREADY,
  m_axi_updates_2_RRESP,
  m_axi_updates_2_RUSER,
  m_axi_updates_2_RVALID,
  m_axi_updates_2_WDATA,
  m_axi_updates_2_WID,
  m_axi_updates_2_WLAST,
  m_axi_updates_2_WREADY,
  m_axi_updates_2_WSTRB,
  m_axi_updates_2_WUSER,
  m_axi_updates_2_WVALID,
  m_axi_updates_3_ARADDR,
  m_axi_updates_3_ARBURST,
  m_axi_updates_3_ARCACHE,
  m_axi_updates_3_ARID,
  m_axi_updates_3_ARLEN,
  m_axi_updates_3_ARLOCK,
  m_axi_updates_3_ARPROT,
  m_axi_updates_3_ARQOS,
  m_axi_updates_3_ARREADY,
  m_axi_updates_3_ARREGION,
  m_axi_updates_3_ARSIZE,
  m_axi_updates_3_ARUSER,
  m_axi_updates_3_ARVALID,
  m_axi_updates_3_AWADDR,
  m_axi_updates_3_AWBURST,
  m_axi_updates_3_AWCACHE,
  m_axi_updates_3_AWID,
  m_axi_updates_3_AWLEN,
  m_axi_updates_3_AWLOCK,
  m_axi_updates_3_AWPROT,
  m_axi_updates_3_AWQOS,
  m_axi_updates_3_AWREADY,
  m_axi_updates_3_AWREGION,
  m_axi_updates_3_AWSIZE,
  m_axi_updates_3_AWUSER,
  m_axi_updates_3_AWVALID,
  m_axi_updates_3_BID,
  m_axi_updates_3_BREADY,
  m_axi_updates_3_BRESP,
  m_axi_updates_3_BUSER,
  m_axi_updates_3_BVALID,
  m_axi_updates_3_RDATA,
  m_axi_updates_3_RID,
  m_axi_updates_3_RLAST,
  m_axi_updates_3_RREADY,
  m_axi_updates_3_RRESP,
  m_axi_updates_3_RUSER,
  m_axi_updates_3_RVALID,
  m_axi_updates_3_WDATA,
  m_axi_updates_3_WID,
  m_axi_updates_3_WLAST,
  m_axi_updates_3_WREADY,
  m_axi_updates_3_WSTRB,
  m_axi_updates_3_WUSER,
  m_axi_updates_3_WVALID,
  m_axi_updates_4_ARADDR,
  m_axi_updates_4_ARBURST,
  m_axi_updates_4_ARCACHE,
  m_axi_updates_4_ARID,
  m_axi_updates_4_ARLEN,
  m_axi_updates_4_ARLOCK,
  m_axi_updates_4_ARPROT,
  m_axi_updates_4_ARQOS,
  m_axi_updates_4_ARREADY,
  m_axi_updates_4_ARREGION,
  m_axi_updates_4_ARSIZE,
  m_axi_updates_4_ARUSER,
  m_axi_updates_4_ARVALID,
  m_axi_updates_4_AWADDR,
  m_axi_updates_4_AWBURST,
  m_axi_updates_4_AWCACHE,
  m_axi_updates_4_AWID,
  m_axi_updates_4_AWLEN,
  m_axi_updates_4_AWLOCK,
  m_axi_updates_4_AWPROT,
  m_axi_updates_4_AWQOS,
  m_axi_updates_4_AWREADY,
  m_axi_updates_4_AWREGION,
  m_axi_updates_4_AWSIZE,
  m_axi_updates_4_AWUSER,
  m_axi_updates_4_AWVALID,
  m_axi_updates_4_BID,
  m_axi_updates_4_BREADY,
  m_axi_updates_4_BRESP,
  m_axi_updates_4_BUSER,
  m_axi_updates_4_BVALID,
  m_axi_updates_4_RDATA,
  m_axi_updates_4_RID,
  m_axi_updates_4_RLAST,
  m_axi_updates_4_RREADY,
  m_axi_updates_4_RRESP,
  m_axi_updates_4_RUSER,
  m_axi_updates_4_RVALID,
  m_axi_updates_4_WDATA,
  m_axi_updates_4_WID,
  m_axi_updates_4_WLAST,
  m_axi_updates_4_WREADY,
  m_axi_updates_4_WSTRB,
  m_axi_updates_4_WUSER,
  m_axi_updates_4_WVALID,
  m_axi_updates_5_ARADDR,
  m_axi_updates_5_ARBURST,
  m_axi_updates_5_ARCACHE,
  m_axi_updates_5_ARID,
  m_axi_updates_5_ARLEN,
  m_axi_updates_5_ARLOCK,
  m_axi_updates_5_ARPROT,
  m_axi_updates_5_ARQOS,
  m_axi_updates_5_ARREADY,
  m_axi_updates_5_ARREGION,
  m_axi_updates_5_ARSIZE,
  m_axi_updates_5_ARUSER,
  m_axi_updates_5_ARVALID,
  m_axi_updates_5_AWADDR,
  m_axi_updates_5_AWBURST,
  m_axi_updates_5_AWCACHE,
  m_axi_updates_5_AWID,
  m_axi_updates_5_AWLEN,
  m_axi_updates_5_AWLOCK,
  m_axi_updates_5_AWPROT,
  m_axi_updates_5_AWQOS,
  m_axi_updates_5_AWREADY,
  m_axi_updates_5_AWREGION,
  m_axi_updates_5_AWSIZE,
  m_axi_updates_5_AWUSER,
  m_axi_updates_5_AWVALID,
  m_axi_updates_5_BID,
  m_axi_updates_5_BREADY,
  m_axi_updates_5_BRESP,
  m_axi_updates_5_BUSER,
  m_axi_updates_5_BVALID,
  m_axi_updates_5_RDATA,
  m_axi_updates_5_RID,
  m_axi_updates_5_RLAST,
  m_axi_updates_5_RREADY,
  m_axi_updates_5_RRESP,
  m_axi_updates_5_RUSER,
  m_axi_updates_5_RVALID,
  m_axi_updates_5_WDATA,
  m_axi_updates_5_WID,
  m_axi_updates_5_WLAST,
  m_axi_updates_5_WREADY,
  m_axi_updates_5_WSTRB,
  m_axi_updates_5_WUSER,
  m_axi_updates_5_WVALID,
  m_axi_updates_6_ARADDR,
  m_axi_updates_6_ARBURST,
  m_axi_updates_6_ARCACHE,
  m_axi_updates_6_ARID,
  m_axi_updates_6_ARLEN,
  m_axi_updates_6_ARLOCK,
  m_axi_updates_6_ARPROT,
  m_axi_updates_6_ARQOS,
  m_axi_updates_6_ARREADY,
  m_axi_updates_6_ARREGION,
  m_axi_updates_6_ARSIZE,
  m_axi_updates_6_ARUSER,
  m_axi_updates_6_ARVALID,
  m_axi_updates_6_AWADDR,
  m_axi_updates_6_AWBURST,
  m_axi_updates_6_AWCACHE,
  m_axi_updates_6_AWID,
  m_axi_updates_6_AWLEN,
  m_axi_updates_6_AWLOCK,
  m_axi_updates_6_AWPROT,
  m_axi_updates_6_AWQOS,
  m_axi_updates_6_AWREADY,
  m_axi_updates_6_AWREGION,
  m_axi_updates_6_AWSIZE,
  m_axi_updates_6_AWUSER,
  m_axi_updates_6_AWVALID,
  m_axi_updates_6_BID,
  m_axi_updates_6_BREADY,
  m_axi_updates_6_BRESP,
  m_axi_updates_6_BUSER,
  m_axi_updates_6_BVALID,
  m_axi_updates_6_RDATA,
  m_axi_updates_6_RID,
  m_axi_updates_6_RLAST,
  m_axi_updates_6_RREADY,
  m_axi_updates_6_RRESP,
  m_axi_updates_6_RUSER,
  m_axi_updates_6_RVALID,
  m_axi_updates_6_WDATA,
  m_axi_updates_6_WID,
  m_axi_updates_6_WLAST,
  m_axi_updates_6_WREADY,
  m_axi_updates_6_WSTRB,
  m_axi_updates_6_WUSER,
  m_axi_updates_6_WVALID,
  m_axi_updates_7_ARADDR,
  m_axi_updates_7_ARBURST,
  m_axi_updates_7_ARCACHE,
  m_axi_updates_7_ARID,
  m_axi_updates_7_ARLEN,
  m_axi_updates_7_ARLOCK,
  m_axi_updates_7_ARPROT,
  m_axi_updates_7_ARQOS,
  m_axi_updates_7_ARREADY,
  m_axi_updates_7_ARREGION,
  m_axi_updates_7_ARSIZE,
  m_axi_updates_7_ARUSER,
  m_axi_updates_7_ARVALID,
  m_axi_updates_7_AWADDR,
  m_axi_updates_7_AWBURST,
  m_axi_updates_7_AWCACHE,
  m_axi_updates_7_AWID,
  m_axi_updates_7_AWLEN,
  m_axi_updates_7_AWLOCK,
  m_axi_updates_7_AWPROT,
  m_axi_updates_7_AWQOS,
  m_axi_updates_7_AWREADY,
  m_axi_updates_7_AWREGION,
  m_axi_updates_7_AWSIZE,
  m_axi_updates_7_AWUSER,
  m_axi_updates_7_AWVALID,
  m_axi_updates_7_BID,
  m_axi_updates_7_BREADY,
  m_axi_updates_7_BRESP,
  m_axi_updates_7_BUSER,
  m_axi_updates_7_BVALID,
  m_axi_updates_7_RDATA,
  m_axi_updates_7_RID,
  m_axi_updates_7_RLAST,
  m_axi_updates_7_RREADY,
  m_axi_updates_7_RRESP,
  m_axi_updates_7_RUSER,
  m_axi_updates_7_RVALID,
  m_axi_updates_7_WDATA,
  m_axi_updates_7_WID,
  m_axi_updates_7_WLAST,
  m_axi_updates_7_WREADY,
  m_axi_updates_7_WSTRB,
  m_axi_updates_7_WUSER,
  m_axi_updates_7_WVALID,
  m_axi_degrees_ARADDR,
  m_axi_degrees_ARBURST,
  m_axi_degrees_ARCACHE,
  m_axi_degrees_ARID,
  m_axi_degrees_ARLEN,
  m_axi_degrees_ARLOCK,
  m_axi_degrees_ARPROT,
  m_axi_degrees_ARQOS,
  m_axi_degrees_ARREADY,
  m_axi_degrees_ARREGION,
  m_axi_degrees_ARSIZE,
  m_axi_degrees_ARUSER,
  m_axi_degrees_ARVALID,
  m_axi_degrees_AWADDR,
  m_axi_degrees_AWBURST,
  m_axi_degrees_AWCACHE,
  m_axi_degrees_AWID,
  m_axi_degrees_AWLEN,
  m_axi_degrees_AWLOCK,
  m_axi_degrees_AWPROT,
  m_axi_degrees_AWQOS,
  m_axi_degrees_AWREADY,
  m_axi_degrees_AWREGION,
  m_axi_degrees_AWSIZE,
  m_axi_degrees_AWUSER,
  m_axi_degrees_AWVALID,
  m_axi_degrees_BID,
  m_axi_degrees_BREADY,
  m_axi_degrees_BRESP,
  m_axi_degrees_BUSER,
  m_axi_degrees_BVALID,
  m_axi_degrees_RDATA,
  m_axi_degrees_RID,
  m_axi_degrees_RLAST,
  m_axi_degrees_RREADY,
  m_axi_degrees_RRESP,
  m_axi_degrees_RUSER,
  m_axi_degrees_RVALID,
  m_axi_degrees_WDATA,
  m_axi_degrees_WID,
  m_axi_degrees_WLAST,
  m_axi_degrees_WREADY,
  m_axi_degrees_WSTRB,
  m_axi_degrees_WUSER,
  m_axi_degrees_WVALID,
  m_axi_rankings_ARADDR,
  m_axi_rankings_ARBURST,
  m_axi_rankings_ARCACHE,
  m_axi_rankings_ARID,
  m_axi_rankings_ARLEN,
  m_axi_rankings_ARLOCK,
  m_axi_rankings_ARPROT,
  m_axi_rankings_ARQOS,
  m_axi_rankings_ARREADY,
  m_axi_rankings_ARREGION,
  m_axi_rankings_ARSIZE,
  m_axi_rankings_ARUSER,
  m_axi_rankings_ARVALID,
  m_axi_rankings_AWADDR,
  m_axi_rankings_AWBURST,
  m_axi_rankings_AWCACHE,
  m_axi_rankings_AWID,
  m_axi_rankings_AWLEN,
  m_axi_rankings_AWLOCK,
  m_axi_rankings_AWPROT,
  m_axi_rankings_AWQOS,
  m_axi_rankings_AWREADY,
  m_axi_rankings_AWREGION,
  m_axi_rankings_AWSIZE,
  m_axi_rankings_AWUSER,
  m_axi_rankings_AWVALID,
  m_axi_rankings_BID,
  m_axi_rankings_BREADY,
  m_axi_rankings_BRESP,
  m_axi_rankings_BUSER,
  m_axi_rankings_BVALID,
  m_axi_rankings_RDATA,
  m_axi_rankings_RID,
  m_axi_rankings_RLAST,
  m_axi_rankings_RREADY,
  m_axi_rankings_RRESP,
  m_axi_rankings_RUSER,
  m_axi_rankings_RVALID,
  m_axi_rankings_WDATA,
  m_axi_rankings_WID,
  m_axi_rankings_WLAST,
  m_axi_rankings_WREADY,
  m_axi_rankings_WSTRB,
  m_axi_rankings_WUSER,
  m_axi_rankings_WVALID,
  m_axi_tmps_ARADDR,
  m_axi_tmps_ARBURST,
  m_axi_tmps_ARCACHE,
  m_axi_tmps_ARID,
  m_axi_tmps_ARLEN,
  m_axi_tmps_ARLOCK,
  m_axi_tmps_ARPROT,
  m_axi_tmps_ARQOS,
  m_axi_tmps_ARREADY,
  m_axi_tmps_ARREGION,
  m_axi_tmps_ARSIZE,
  m_axi_tmps_ARUSER,
  m_axi_tmps_ARVALID,
  m_axi_tmps_AWADDR,
  m_axi_tmps_AWBURST,
  m_axi_tmps_AWCACHE,
  m_axi_tmps_AWID,
  m_axi_tmps_AWLEN,
  m_axi_tmps_AWLOCK,
  m_axi_tmps_AWPROT,
  m_axi_tmps_AWQOS,
  m_axi_tmps_AWREADY,
  m_axi_tmps_AWREGION,
  m_axi_tmps_AWSIZE,
  m_axi_tmps_AWUSER,
  m_axi_tmps_AWVALID,
  m_axi_tmps_BID,
  m_axi_tmps_BREADY,
  m_axi_tmps_BRESP,
  m_axi_tmps_BUSER,
  m_axi_tmps_BVALID,
  m_axi_tmps_RDATA,
  m_axi_tmps_RID,
  m_axi_tmps_RLAST,
  m_axi_tmps_RREADY,
  m_axi_tmps_RRESP,
  m_axi_tmps_RUSER,
  m_axi_tmps_RVALID,
  m_axi_tmps_WDATA,
  m_axi_tmps_WID,
  m_axi_tmps_WLAST,
  m_axi_tmps_WREADY,
  m_axi_tmps_WSTRB,
  m_axi_tmps_WUSER,
  m_axi_tmps_WVALID
);

  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 9;
  parameter C_S_AXI_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
  parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
  input ap_clk;
  input ap_rst_n;
  input s_axi_control_AWVALID;
  output s_axi_control_AWREADY;
  input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_AWADDR;
  input s_axi_control_WVALID;
  output s_axi_control_WREADY;
  input [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_WDATA;
  input [C_S_AXI_CONTROL_WSTRB_WIDTH-1:0] s_axi_control_WSTRB;
  input s_axi_control_ARVALID;
  output s_axi_control_ARREADY;
  input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_ARADDR;
  output s_axi_control_RVALID;
  input s_axi_control_RREADY;
  output [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_RDATA;
  output [1:0] s_axi_control_RRESP;
  output s_axi_control_BVALID;
  input s_axi_control_BREADY;
  output [1:0] s_axi_control_BRESP;
  output interrupt;
  output [63:0] m_axi_metadata_ARADDR;
  output [1:0] m_axi_metadata_ARBURST;
  output [3:0] m_axi_metadata_ARCACHE;
  output [0:0] m_axi_metadata_ARID;
  output [7:0] m_axi_metadata_ARLEN;
  output m_axi_metadata_ARLOCK;
  output [2:0] m_axi_metadata_ARPROT;
  output [3:0] m_axi_metadata_ARQOS;
  input m_axi_metadata_ARREADY;
  output [3:0] m_axi_metadata_ARREGION;
  output [2:0] m_axi_metadata_ARSIZE;
  output m_axi_metadata_ARUSER;
  output m_axi_metadata_ARVALID;
  output [63:0] m_axi_metadata_AWADDR;
  output [1:0] m_axi_metadata_AWBURST;
  output [3:0] m_axi_metadata_AWCACHE;
  output [0:0] m_axi_metadata_AWID;
  output [7:0] m_axi_metadata_AWLEN;
  output m_axi_metadata_AWLOCK;
  output [2:0] m_axi_metadata_AWPROT;
  output [3:0] m_axi_metadata_AWQOS;
  input m_axi_metadata_AWREADY;
  output [3:0] m_axi_metadata_AWREGION;
  output [2:0] m_axi_metadata_AWSIZE;
  output m_axi_metadata_AWUSER;
  output m_axi_metadata_AWVALID;
  input [0:0] m_axi_metadata_BID;
  output m_axi_metadata_BREADY;
  input [1:0] m_axi_metadata_BRESP;
  input m_axi_metadata_BUSER;
  input m_axi_metadata_BVALID;
  input [63:0] m_axi_metadata_RDATA;
  input [0:0] m_axi_metadata_RID;
  input m_axi_metadata_RLAST;
  output m_axi_metadata_RREADY;
  input [1:0] m_axi_metadata_RRESP;
  input m_axi_metadata_RUSER;
  input m_axi_metadata_RVALID;
  output [63:0] m_axi_metadata_WDATA;
  output [0:0] m_axi_metadata_WID;
  output m_axi_metadata_WLAST;
  input m_axi_metadata_WREADY;
  output [7:0] m_axi_metadata_WSTRB;
  output m_axi_metadata_WUSER;
  output m_axi_metadata_WVALID;
  output [63:0] m_axi_edges_0_ARADDR;
  output [1:0] m_axi_edges_0_ARBURST;
  output [3:0] m_axi_edges_0_ARCACHE;
  output [0:0] m_axi_edges_0_ARID;
  output [7:0] m_axi_edges_0_ARLEN;
  output m_axi_edges_0_ARLOCK;
  output [2:0] m_axi_edges_0_ARPROT;
  output [3:0] m_axi_edges_0_ARQOS;
  input m_axi_edges_0_ARREADY;
  output [3:0] m_axi_edges_0_ARREGION;
  output [2:0] m_axi_edges_0_ARSIZE;
  output m_axi_edges_0_ARUSER;
  output m_axi_edges_0_ARVALID;
  output [63:0] m_axi_edges_0_AWADDR;
  output [1:0] m_axi_edges_0_AWBURST;
  output [3:0] m_axi_edges_0_AWCACHE;
  output [0:0] m_axi_edges_0_AWID;
  output [7:0] m_axi_edges_0_AWLEN;
  output m_axi_edges_0_AWLOCK;
  output [2:0] m_axi_edges_0_AWPROT;
  output [3:0] m_axi_edges_0_AWQOS;
  input m_axi_edges_0_AWREADY;
  output [3:0] m_axi_edges_0_AWREGION;
  output [2:0] m_axi_edges_0_AWSIZE;
  output m_axi_edges_0_AWUSER;
  output m_axi_edges_0_AWVALID;
  input [0:0] m_axi_edges_0_BID;
  output m_axi_edges_0_BREADY;
  input [1:0] m_axi_edges_0_BRESP;
  input m_axi_edges_0_BUSER;
  input m_axi_edges_0_BVALID;
  input [511:0] m_axi_edges_0_RDATA;
  input [0:0] m_axi_edges_0_RID;
  input m_axi_edges_0_RLAST;
  output m_axi_edges_0_RREADY;
  input [1:0] m_axi_edges_0_RRESP;
  input m_axi_edges_0_RUSER;
  input m_axi_edges_0_RVALID;
  output [511:0] m_axi_edges_0_WDATA;
  output [0:0] m_axi_edges_0_WID;
  output m_axi_edges_0_WLAST;
  input m_axi_edges_0_WREADY;
  output [63:0] m_axi_edges_0_WSTRB;
  output m_axi_edges_0_WUSER;
  output m_axi_edges_0_WVALID;
  output [63:0] m_axi_edges_1_ARADDR;
  output [1:0] m_axi_edges_1_ARBURST;
  output [3:0] m_axi_edges_1_ARCACHE;
  output [0:0] m_axi_edges_1_ARID;
  output [7:0] m_axi_edges_1_ARLEN;
  output m_axi_edges_1_ARLOCK;
  output [2:0] m_axi_edges_1_ARPROT;
  output [3:0] m_axi_edges_1_ARQOS;
  input m_axi_edges_1_ARREADY;
  output [3:0] m_axi_edges_1_ARREGION;
  output [2:0] m_axi_edges_1_ARSIZE;
  output m_axi_edges_1_ARUSER;
  output m_axi_edges_1_ARVALID;
  output [63:0] m_axi_edges_1_AWADDR;
  output [1:0] m_axi_edges_1_AWBURST;
  output [3:0] m_axi_edges_1_AWCACHE;
  output [0:0] m_axi_edges_1_AWID;
  output [7:0] m_axi_edges_1_AWLEN;
  output m_axi_edges_1_AWLOCK;
  output [2:0] m_axi_edges_1_AWPROT;
  output [3:0] m_axi_edges_1_AWQOS;
  input m_axi_edges_1_AWREADY;
  output [3:0] m_axi_edges_1_AWREGION;
  output [2:0] m_axi_edges_1_AWSIZE;
  output m_axi_edges_1_AWUSER;
  output m_axi_edges_1_AWVALID;
  input [0:0] m_axi_edges_1_BID;
  output m_axi_edges_1_BREADY;
  input [1:0] m_axi_edges_1_BRESP;
  input m_axi_edges_1_BUSER;
  input m_axi_edges_1_BVALID;
  input [511:0] m_axi_edges_1_RDATA;
  input [0:0] m_axi_edges_1_RID;
  input m_axi_edges_1_RLAST;
  output m_axi_edges_1_RREADY;
  input [1:0] m_axi_edges_1_RRESP;
  input m_axi_edges_1_RUSER;
  input m_axi_edges_1_RVALID;
  output [511:0] m_axi_edges_1_WDATA;
  output [0:0] m_axi_edges_1_WID;
  output m_axi_edges_1_WLAST;
  input m_axi_edges_1_WREADY;
  output [63:0] m_axi_edges_1_WSTRB;
  output m_axi_edges_1_WUSER;
  output m_axi_edges_1_WVALID;
  output [63:0] m_axi_edges_2_ARADDR;
  output [1:0] m_axi_edges_2_ARBURST;
  output [3:0] m_axi_edges_2_ARCACHE;
  output [0:0] m_axi_edges_2_ARID;
  output [7:0] m_axi_edges_2_ARLEN;
  output m_axi_edges_2_ARLOCK;
  output [2:0] m_axi_edges_2_ARPROT;
  output [3:0] m_axi_edges_2_ARQOS;
  input m_axi_edges_2_ARREADY;
  output [3:0] m_axi_edges_2_ARREGION;
  output [2:0] m_axi_edges_2_ARSIZE;
  output m_axi_edges_2_ARUSER;
  output m_axi_edges_2_ARVALID;
  output [63:0] m_axi_edges_2_AWADDR;
  output [1:0] m_axi_edges_2_AWBURST;
  output [3:0] m_axi_edges_2_AWCACHE;
  output [0:0] m_axi_edges_2_AWID;
  output [7:0] m_axi_edges_2_AWLEN;
  output m_axi_edges_2_AWLOCK;
  output [2:0] m_axi_edges_2_AWPROT;
  output [3:0] m_axi_edges_2_AWQOS;
  input m_axi_edges_2_AWREADY;
  output [3:0] m_axi_edges_2_AWREGION;
  output [2:0] m_axi_edges_2_AWSIZE;
  output m_axi_edges_2_AWUSER;
  output m_axi_edges_2_AWVALID;
  input [0:0] m_axi_edges_2_BID;
  output m_axi_edges_2_BREADY;
  input [1:0] m_axi_edges_2_BRESP;
  input m_axi_edges_2_BUSER;
  input m_axi_edges_2_BVALID;
  input [511:0] m_axi_edges_2_RDATA;
  input [0:0] m_axi_edges_2_RID;
  input m_axi_edges_2_RLAST;
  output m_axi_edges_2_RREADY;
  input [1:0] m_axi_edges_2_RRESP;
  input m_axi_edges_2_RUSER;
  input m_axi_edges_2_RVALID;
  output [511:0] m_axi_edges_2_WDATA;
  output [0:0] m_axi_edges_2_WID;
  output m_axi_edges_2_WLAST;
  input m_axi_edges_2_WREADY;
  output [63:0] m_axi_edges_2_WSTRB;
  output m_axi_edges_2_WUSER;
  output m_axi_edges_2_WVALID;
  output [63:0] m_axi_edges_3_ARADDR;
  output [1:0] m_axi_edges_3_ARBURST;
  output [3:0] m_axi_edges_3_ARCACHE;
  output [0:0] m_axi_edges_3_ARID;
  output [7:0] m_axi_edges_3_ARLEN;
  output m_axi_edges_3_ARLOCK;
  output [2:0] m_axi_edges_3_ARPROT;
  output [3:0] m_axi_edges_3_ARQOS;
  input m_axi_edges_3_ARREADY;
  output [3:0] m_axi_edges_3_ARREGION;
  output [2:0] m_axi_edges_3_ARSIZE;
  output m_axi_edges_3_ARUSER;
  output m_axi_edges_3_ARVALID;
  output [63:0] m_axi_edges_3_AWADDR;
  output [1:0] m_axi_edges_3_AWBURST;
  output [3:0] m_axi_edges_3_AWCACHE;
  output [0:0] m_axi_edges_3_AWID;
  output [7:0] m_axi_edges_3_AWLEN;
  output m_axi_edges_3_AWLOCK;
  output [2:0] m_axi_edges_3_AWPROT;
  output [3:0] m_axi_edges_3_AWQOS;
  input m_axi_edges_3_AWREADY;
  output [3:0] m_axi_edges_3_AWREGION;
  output [2:0] m_axi_edges_3_AWSIZE;
  output m_axi_edges_3_AWUSER;
  output m_axi_edges_3_AWVALID;
  input [0:0] m_axi_edges_3_BID;
  output m_axi_edges_3_BREADY;
  input [1:0] m_axi_edges_3_BRESP;
  input m_axi_edges_3_BUSER;
  input m_axi_edges_3_BVALID;
  input [511:0] m_axi_edges_3_RDATA;
  input [0:0] m_axi_edges_3_RID;
  input m_axi_edges_3_RLAST;
  output m_axi_edges_3_RREADY;
  input [1:0] m_axi_edges_3_RRESP;
  input m_axi_edges_3_RUSER;
  input m_axi_edges_3_RVALID;
  output [511:0] m_axi_edges_3_WDATA;
  output [0:0] m_axi_edges_3_WID;
  output m_axi_edges_3_WLAST;
  input m_axi_edges_3_WREADY;
  output [63:0] m_axi_edges_3_WSTRB;
  output m_axi_edges_3_WUSER;
  output m_axi_edges_3_WVALID;
  output [63:0] m_axi_edges_4_ARADDR;
  output [1:0] m_axi_edges_4_ARBURST;
  output [3:0] m_axi_edges_4_ARCACHE;
  output [0:0] m_axi_edges_4_ARID;
  output [7:0] m_axi_edges_4_ARLEN;
  output m_axi_edges_4_ARLOCK;
  output [2:0] m_axi_edges_4_ARPROT;
  output [3:0] m_axi_edges_4_ARQOS;
  input m_axi_edges_4_ARREADY;
  output [3:0] m_axi_edges_4_ARREGION;
  output [2:0] m_axi_edges_4_ARSIZE;
  output m_axi_edges_4_ARUSER;
  output m_axi_edges_4_ARVALID;
  output [63:0] m_axi_edges_4_AWADDR;
  output [1:0] m_axi_edges_4_AWBURST;
  output [3:0] m_axi_edges_4_AWCACHE;
  output [0:0] m_axi_edges_4_AWID;
  output [7:0] m_axi_edges_4_AWLEN;
  output m_axi_edges_4_AWLOCK;
  output [2:0] m_axi_edges_4_AWPROT;
  output [3:0] m_axi_edges_4_AWQOS;
  input m_axi_edges_4_AWREADY;
  output [3:0] m_axi_edges_4_AWREGION;
  output [2:0] m_axi_edges_4_AWSIZE;
  output m_axi_edges_4_AWUSER;
  output m_axi_edges_4_AWVALID;
  input [0:0] m_axi_edges_4_BID;
  output m_axi_edges_4_BREADY;
  input [1:0] m_axi_edges_4_BRESP;
  input m_axi_edges_4_BUSER;
  input m_axi_edges_4_BVALID;
  input [511:0] m_axi_edges_4_RDATA;
  input [0:0] m_axi_edges_4_RID;
  input m_axi_edges_4_RLAST;
  output m_axi_edges_4_RREADY;
  input [1:0] m_axi_edges_4_RRESP;
  input m_axi_edges_4_RUSER;
  input m_axi_edges_4_RVALID;
  output [511:0] m_axi_edges_4_WDATA;
  output [0:0] m_axi_edges_4_WID;
  output m_axi_edges_4_WLAST;
  input m_axi_edges_4_WREADY;
  output [63:0] m_axi_edges_4_WSTRB;
  output m_axi_edges_4_WUSER;
  output m_axi_edges_4_WVALID;
  output [63:0] m_axi_edges_5_ARADDR;
  output [1:0] m_axi_edges_5_ARBURST;
  output [3:0] m_axi_edges_5_ARCACHE;
  output [0:0] m_axi_edges_5_ARID;
  output [7:0] m_axi_edges_5_ARLEN;
  output m_axi_edges_5_ARLOCK;
  output [2:0] m_axi_edges_5_ARPROT;
  output [3:0] m_axi_edges_5_ARQOS;
  input m_axi_edges_5_ARREADY;
  output [3:0] m_axi_edges_5_ARREGION;
  output [2:0] m_axi_edges_5_ARSIZE;
  output m_axi_edges_5_ARUSER;
  output m_axi_edges_5_ARVALID;
  output [63:0] m_axi_edges_5_AWADDR;
  output [1:0] m_axi_edges_5_AWBURST;
  output [3:0] m_axi_edges_5_AWCACHE;
  output [0:0] m_axi_edges_5_AWID;
  output [7:0] m_axi_edges_5_AWLEN;
  output m_axi_edges_5_AWLOCK;
  output [2:0] m_axi_edges_5_AWPROT;
  output [3:0] m_axi_edges_5_AWQOS;
  input m_axi_edges_5_AWREADY;
  output [3:0] m_axi_edges_5_AWREGION;
  output [2:0] m_axi_edges_5_AWSIZE;
  output m_axi_edges_5_AWUSER;
  output m_axi_edges_5_AWVALID;
  input [0:0] m_axi_edges_5_BID;
  output m_axi_edges_5_BREADY;
  input [1:0] m_axi_edges_5_BRESP;
  input m_axi_edges_5_BUSER;
  input m_axi_edges_5_BVALID;
  input [511:0] m_axi_edges_5_RDATA;
  input [0:0] m_axi_edges_5_RID;
  input m_axi_edges_5_RLAST;
  output m_axi_edges_5_RREADY;
  input [1:0] m_axi_edges_5_RRESP;
  input m_axi_edges_5_RUSER;
  input m_axi_edges_5_RVALID;
  output [511:0] m_axi_edges_5_WDATA;
  output [0:0] m_axi_edges_5_WID;
  output m_axi_edges_5_WLAST;
  input m_axi_edges_5_WREADY;
  output [63:0] m_axi_edges_5_WSTRB;
  output m_axi_edges_5_WUSER;
  output m_axi_edges_5_WVALID;
  output [63:0] m_axi_edges_6_ARADDR;
  output [1:0] m_axi_edges_6_ARBURST;
  output [3:0] m_axi_edges_6_ARCACHE;
  output [0:0] m_axi_edges_6_ARID;
  output [7:0] m_axi_edges_6_ARLEN;
  output m_axi_edges_6_ARLOCK;
  output [2:0] m_axi_edges_6_ARPROT;
  output [3:0] m_axi_edges_6_ARQOS;
  input m_axi_edges_6_ARREADY;
  output [3:0] m_axi_edges_6_ARREGION;
  output [2:0] m_axi_edges_6_ARSIZE;
  output m_axi_edges_6_ARUSER;
  output m_axi_edges_6_ARVALID;
  output [63:0] m_axi_edges_6_AWADDR;
  output [1:0] m_axi_edges_6_AWBURST;
  output [3:0] m_axi_edges_6_AWCACHE;
  output [0:0] m_axi_edges_6_AWID;
  output [7:0] m_axi_edges_6_AWLEN;
  output m_axi_edges_6_AWLOCK;
  output [2:0] m_axi_edges_6_AWPROT;
  output [3:0] m_axi_edges_6_AWQOS;
  input m_axi_edges_6_AWREADY;
  output [3:0] m_axi_edges_6_AWREGION;
  output [2:0] m_axi_edges_6_AWSIZE;
  output m_axi_edges_6_AWUSER;
  output m_axi_edges_6_AWVALID;
  input [0:0] m_axi_edges_6_BID;
  output m_axi_edges_6_BREADY;
  input [1:0] m_axi_edges_6_BRESP;
  input m_axi_edges_6_BUSER;
  input m_axi_edges_6_BVALID;
  input [511:0] m_axi_edges_6_RDATA;
  input [0:0] m_axi_edges_6_RID;
  input m_axi_edges_6_RLAST;
  output m_axi_edges_6_RREADY;
  input [1:0] m_axi_edges_6_RRESP;
  input m_axi_edges_6_RUSER;
  input m_axi_edges_6_RVALID;
  output [511:0] m_axi_edges_6_WDATA;
  output [0:0] m_axi_edges_6_WID;
  output m_axi_edges_6_WLAST;
  input m_axi_edges_6_WREADY;
  output [63:0] m_axi_edges_6_WSTRB;
  output m_axi_edges_6_WUSER;
  output m_axi_edges_6_WVALID;
  output [63:0] m_axi_edges_7_ARADDR;
  output [1:0] m_axi_edges_7_ARBURST;
  output [3:0] m_axi_edges_7_ARCACHE;
  output [0:0] m_axi_edges_7_ARID;
  output [7:0] m_axi_edges_7_ARLEN;
  output m_axi_edges_7_ARLOCK;
  output [2:0] m_axi_edges_7_ARPROT;
  output [3:0] m_axi_edges_7_ARQOS;
  input m_axi_edges_7_ARREADY;
  output [3:0] m_axi_edges_7_ARREGION;
  output [2:0] m_axi_edges_7_ARSIZE;
  output m_axi_edges_7_ARUSER;
  output m_axi_edges_7_ARVALID;
  output [63:0] m_axi_edges_7_AWADDR;
  output [1:0] m_axi_edges_7_AWBURST;
  output [3:0] m_axi_edges_7_AWCACHE;
  output [0:0] m_axi_edges_7_AWID;
  output [7:0] m_axi_edges_7_AWLEN;
  output m_axi_edges_7_AWLOCK;
  output [2:0] m_axi_edges_7_AWPROT;
  output [3:0] m_axi_edges_7_AWQOS;
  input m_axi_edges_7_AWREADY;
  output [3:0] m_axi_edges_7_AWREGION;
  output [2:0] m_axi_edges_7_AWSIZE;
  output m_axi_edges_7_AWUSER;
  output m_axi_edges_7_AWVALID;
  input [0:0] m_axi_edges_7_BID;
  output m_axi_edges_7_BREADY;
  input [1:0] m_axi_edges_7_BRESP;
  input m_axi_edges_7_BUSER;
  input m_axi_edges_7_BVALID;
  input [511:0] m_axi_edges_7_RDATA;
  input [0:0] m_axi_edges_7_RID;
  input m_axi_edges_7_RLAST;
  output m_axi_edges_7_RREADY;
  input [1:0] m_axi_edges_7_RRESP;
  input m_axi_edges_7_RUSER;
  input m_axi_edges_7_RVALID;
  output [511:0] m_axi_edges_7_WDATA;
  output [0:0] m_axi_edges_7_WID;
  output m_axi_edges_7_WLAST;
  input m_axi_edges_7_WREADY;
  output [63:0] m_axi_edges_7_WSTRB;
  output m_axi_edges_7_WUSER;
  output m_axi_edges_7_WVALID;
  output [63:0] m_axi_updates_0_ARADDR;
  output [1:0] m_axi_updates_0_ARBURST;
  output [3:0] m_axi_updates_0_ARCACHE;
  output [0:0] m_axi_updates_0_ARID;
  output [7:0] m_axi_updates_0_ARLEN;
  output m_axi_updates_0_ARLOCK;
  output [2:0] m_axi_updates_0_ARPROT;
  output [3:0] m_axi_updates_0_ARQOS;
  input m_axi_updates_0_ARREADY;
  output [3:0] m_axi_updates_0_ARREGION;
  output [2:0] m_axi_updates_0_ARSIZE;
  output m_axi_updates_0_ARUSER;
  output m_axi_updates_0_ARVALID;
  output [63:0] m_axi_updates_0_AWADDR;
  output [1:0] m_axi_updates_0_AWBURST;
  output [3:0] m_axi_updates_0_AWCACHE;
  output [0:0] m_axi_updates_0_AWID;
  output [7:0] m_axi_updates_0_AWLEN;
  output m_axi_updates_0_AWLOCK;
  output [2:0] m_axi_updates_0_AWPROT;
  output [3:0] m_axi_updates_0_AWQOS;
  input m_axi_updates_0_AWREADY;
  output [3:0] m_axi_updates_0_AWREGION;
  output [2:0] m_axi_updates_0_AWSIZE;
  output m_axi_updates_0_AWUSER;
  output m_axi_updates_0_AWVALID;
  input [0:0] m_axi_updates_0_BID;
  output m_axi_updates_0_BREADY;
  input [1:0] m_axi_updates_0_BRESP;
  input m_axi_updates_0_BUSER;
  input m_axi_updates_0_BVALID;
  input [511:0] m_axi_updates_0_RDATA;
  input [0:0] m_axi_updates_0_RID;
  input m_axi_updates_0_RLAST;
  output m_axi_updates_0_RREADY;
  input [1:0] m_axi_updates_0_RRESP;
  input m_axi_updates_0_RUSER;
  input m_axi_updates_0_RVALID;
  output [511:0] m_axi_updates_0_WDATA;
  output [0:0] m_axi_updates_0_WID;
  output m_axi_updates_0_WLAST;
  input m_axi_updates_0_WREADY;
  output [63:0] m_axi_updates_0_WSTRB;
  output m_axi_updates_0_WUSER;
  output m_axi_updates_0_WVALID;
  output [63:0] m_axi_updates_1_ARADDR;
  output [1:0] m_axi_updates_1_ARBURST;
  output [3:0] m_axi_updates_1_ARCACHE;
  output [0:0] m_axi_updates_1_ARID;
  output [7:0] m_axi_updates_1_ARLEN;
  output m_axi_updates_1_ARLOCK;
  output [2:0] m_axi_updates_1_ARPROT;
  output [3:0] m_axi_updates_1_ARQOS;
  input m_axi_updates_1_ARREADY;
  output [3:0] m_axi_updates_1_ARREGION;
  output [2:0] m_axi_updates_1_ARSIZE;
  output m_axi_updates_1_ARUSER;
  output m_axi_updates_1_ARVALID;
  output [63:0] m_axi_updates_1_AWADDR;
  output [1:0] m_axi_updates_1_AWBURST;
  output [3:0] m_axi_updates_1_AWCACHE;
  output [0:0] m_axi_updates_1_AWID;
  output [7:0] m_axi_updates_1_AWLEN;
  output m_axi_updates_1_AWLOCK;
  output [2:0] m_axi_updates_1_AWPROT;
  output [3:0] m_axi_updates_1_AWQOS;
  input m_axi_updates_1_AWREADY;
  output [3:0] m_axi_updates_1_AWREGION;
  output [2:0] m_axi_updates_1_AWSIZE;
  output m_axi_updates_1_AWUSER;
  output m_axi_updates_1_AWVALID;
  input [0:0] m_axi_updates_1_BID;
  output m_axi_updates_1_BREADY;
  input [1:0] m_axi_updates_1_BRESP;
  input m_axi_updates_1_BUSER;
  input m_axi_updates_1_BVALID;
  input [511:0] m_axi_updates_1_RDATA;
  input [0:0] m_axi_updates_1_RID;
  input m_axi_updates_1_RLAST;
  output m_axi_updates_1_RREADY;
  input [1:0] m_axi_updates_1_RRESP;
  input m_axi_updates_1_RUSER;
  input m_axi_updates_1_RVALID;
  output [511:0] m_axi_updates_1_WDATA;
  output [0:0] m_axi_updates_1_WID;
  output m_axi_updates_1_WLAST;
  input m_axi_updates_1_WREADY;
  output [63:0] m_axi_updates_1_WSTRB;
  output m_axi_updates_1_WUSER;
  output m_axi_updates_1_WVALID;
  output [63:0] m_axi_updates_2_ARADDR;
  output [1:0] m_axi_updates_2_ARBURST;
  output [3:0] m_axi_updates_2_ARCACHE;
  output [0:0] m_axi_updates_2_ARID;
  output [7:0] m_axi_updates_2_ARLEN;
  output m_axi_updates_2_ARLOCK;
  output [2:0] m_axi_updates_2_ARPROT;
  output [3:0] m_axi_updates_2_ARQOS;
  input m_axi_updates_2_ARREADY;
  output [3:0] m_axi_updates_2_ARREGION;
  output [2:0] m_axi_updates_2_ARSIZE;
  output m_axi_updates_2_ARUSER;
  output m_axi_updates_2_ARVALID;
  output [63:0] m_axi_updates_2_AWADDR;
  output [1:0] m_axi_updates_2_AWBURST;
  output [3:0] m_axi_updates_2_AWCACHE;
  output [0:0] m_axi_updates_2_AWID;
  output [7:0] m_axi_updates_2_AWLEN;
  output m_axi_updates_2_AWLOCK;
  output [2:0] m_axi_updates_2_AWPROT;
  output [3:0] m_axi_updates_2_AWQOS;
  input m_axi_updates_2_AWREADY;
  output [3:0] m_axi_updates_2_AWREGION;
  output [2:0] m_axi_updates_2_AWSIZE;
  output m_axi_updates_2_AWUSER;
  output m_axi_updates_2_AWVALID;
  input [0:0] m_axi_updates_2_BID;
  output m_axi_updates_2_BREADY;
  input [1:0] m_axi_updates_2_BRESP;
  input m_axi_updates_2_BUSER;
  input m_axi_updates_2_BVALID;
  input [511:0] m_axi_updates_2_RDATA;
  input [0:0] m_axi_updates_2_RID;
  input m_axi_updates_2_RLAST;
  output m_axi_updates_2_RREADY;
  input [1:0] m_axi_updates_2_RRESP;
  input m_axi_updates_2_RUSER;
  input m_axi_updates_2_RVALID;
  output [511:0] m_axi_updates_2_WDATA;
  output [0:0] m_axi_updates_2_WID;
  output m_axi_updates_2_WLAST;
  input m_axi_updates_2_WREADY;
  output [63:0] m_axi_updates_2_WSTRB;
  output m_axi_updates_2_WUSER;
  output m_axi_updates_2_WVALID;
  output [63:0] m_axi_updates_3_ARADDR;
  output [1:0] m_axi_updates_3_ARBURST;
  output [3:0] m_axi_updates_3_ARCACHE;
  output [0:0] m_axi_updates_3_ARID;
  output [7:0] m_axi_updates_3_ARLEN;
  output m_axi_updates_3_ARLOCK;
  output [2:0] m_axi_updates_3_ARPROT;
  output [3:0] m_axi_updates_3_ARQOS;
  input m_axi_updates_3_ARREADY;
  output [3:0] m_axi_updates_3_ARREGION;
  output [2:0] m_axi_updates_3_ARSIZE;
  output m_axi_updates_3_ARUSER;
  output m_axi_updates_3_ARVALID;
  output [63:0] m_axi_updates_3_AWADDR;
  output [1:0] m_axi_updates_3_AWBURST;
  output [3:0] m_axi_updates_3_AWCACHE;
  output [0:0] m_axi_updates_3_AWID;
  output [7:0] m_axi_updates_3_AWLEN;
  output m_axi_updates_3_AWLOCK;
  output [2:0] m_axi_updates_3_AWPROT;
  output [3:0] m_axi_updates_3_AWQOS;
  input m_axi_updates_3_AWREADY;
  output [3:0] m_axi_updates_3_AWREGION;
  output [2:0] m_axi_updates_3_AWSIZE;
  output m_axi_updates_3_AWUSER;
  output m_axi_updates_3_AWVALID;
  input [0:0] m_axi_updates_3_BID;
  output m_axi_updates_3_BREADY;
  input [1:0] m_axi_updates_3_BRESP;
  input m_axi_updates_3_BUSER;
  input m_axi_updates_3_BVALID;
  input [511:0] m_axi_updates_3_RDATA;
  input [0:0] m_axi_updates_3_RID;
  input m_axi_updates_3_RLAST;
  output m_axi_updates_3_RREADY;
  input [1:0] m_axi_updates_3_RRESP;
  input m_axi_updates_3_RUSER;
  input m_axi_updates_3_RVALID;
  output [511:0] m_axi_updates_3_WDATA;
  output [0:0] m_axi_updates_3_WID;
  output m_axi_updates_3_WLAST;
  input m_axi_updates_3_WREADY;
  output [63:0] m_axi_updates_3_WSTRB;
  output m_axi_updates_3_WUSER;
  output m_axi_updates_3_WVALID;
  output [63:0] m_axi_updates_4_ARADDR;
  output [1:0] m_axi_updates_4_ARBURST;
  output [3:0] m_axi_updates_4_ARCACHE;
  output [0:0] m_axi_updates_4_ARID;
  output [7:0] m_axi_updates_4_ARLEN;
  output m_axi_updates_4_ARLOCK;
  output [2:0] m_axi_updates_4_ARPROT;
  output [3:0] m_axi_updates_4_ARQOS;
  input m_axi_updates_4_ARREADY;
  output [3:0] m_axi_updates_4_ARREGION;
  output [2:0] m_axi_updates_4_ARSIZE;
  output m_axi_updates_4_ARUSER;
  output m_axi_updates_4_ARVALID;
  output [63:0] m_axi_updates_4_AWADDR;
  output [1:0] m_axi_updates_4_AWBURST;
  output [3:0] m_axi_updates_4_AWCACHE;
  output [0:0] m_axi_updates_4_AWID;
  output [7:0] m_axi_updates_4_AWLEN;
  output m_axi_updates_4_AWLOCK;
  output [2:0] m_axi_updates_4_AWPROT;
  output [3:0] m_axi_updates_4_AWQOS;
  input m_axi_updates_4_AWREADY;
  output [3:0] m_axi_updates_4_AWREGION;
  output [2:0] m_axi_updates_4_AWSIZE;
  output m_axi_updates_4_AWUSER;
  output m_axi_updates_4_AWVALID;
  input [0:0] m_axi_updates_4_BID;
  output m_axi_updates_4_BREADY;
  input [1:0] m_axi_updates_4_BRESP;
  input m_axi_updates_4_BUSER;
  input m_axi_updates_4_BVALID;
  input [511:0] m_axi_updates_4_RDATA;
  input [0:0] m_axi_updates_4_RID;
  input m_axi_updates_4_RLAST;
  output m_axi_updates_4_RREADY;
  input [1:0] m_axi_updates_4_RRESP;
  input m_axi_updates_4_RUSER;
  input m_axi_updates_4_RVALID;
  output [511:0] m_axi_updates_4_WDATA;
  output [0:0] m_axi_updates_4_WID;
  output m_axi_updates_4_WLAST;
  input m_axi_updates_4_WREADY;
  output [63:0] m_axi_updates_4_WSTRB;
  output m_axi_updates_4_WUSER;
  output m_axi_updates_4_WVALID;
  output [63:0] m_axi_updates_5_ARADDR;
  output [1:0] m_axi_updates_5_ARBURST;
  output [3:0] m_axi_updates_5_ARCACHE;
  output [0:0] m_axi_updates_5_ARID;
  output [7:0] m_axi_updates_5_ARLEN;
  output m_axi_updates_5_ARLOCK;
  output [2:0] m_axi_updates_5_ARPROT;
  output [3:0] m_axi_updates_5_ARQOS;
  input m_axi_updates_5_ARREADY;
  output [3:0] m_axi_updates_5_ARREGION;
  output [2:0] m_axi_updates_5_ARSIZE;
  output m_axi_updates_5_ARUSER;
  output m_axi_updates_5_ARVALID;
  output [63:0] m_axi_updates_5_AWADDR;
  output [1:0] m_axi_updates_5_AWBURST;
  output [3:0] m_axi_updates_5_AWCACHE;
  output [0:0] m_axi_updates_5_AWID;
  output [7:0] m_axi_updates_5_AWLEN;
  output m_axi_updates_5_AWLOCK;
  output [2:0] m_axi_updates_5_AWPROT;
  output [3:0] m_axi_updates_5_AWQOS;
  input m_axi_updates_5_AWREADY;
  output [3:0] m_axi_updates_5_AWREGION;
  output [2:0] m_axi_updates_5_AWSIZE;
  output m_axi_updates_5_AWUSER;
  output m_axi_updates_5_AWVALID;
  input [0:0] m_axi_updates_5_BID;
  output m_axi_updates_5_BREADY;
  input [1:0] m_axi_updates_5_BRESP;
  input m_axi_updates_5_BUSER;
  input m_axi_updates_5_BVALID;
  input [511:0] m_axi_updates_5_RDATA;
  input [0:0] m_axi_updates_5_RID;
  input m_axi_updates_5_RLAST;
  output m_axi_updates_5_RREADY;
  input [1:0] m_axi_updates_5_RRESP;
  input m_axi_updates_5_RUSER;
  input m_axi_updates_5_RVALID;
  output [511:0] m_axi_updates_5_WDATA;
  output [0:0] m_axi_updates_5_WID;
  output m_axi_updates_5_WLAST;
  input m_axi_updates_5_WREADY;
  output [63:0] m_axi_updates_5_WSTRB;
  output m_axi_updates_5_WUSER;
  output m_axi_updates_5_WVALID;
  output [63:0] m_axi_updates_6_ARADDR;
  output [1:0] m_axi_updates_6_ARBURST;
  output [3:0] m_axi_updates_6_ARCACHE;
  output [0:0] m_axi_updates_6_ARID;
  output [7:0] m_axi_updates_6_ARLEN;
  output m_axi_updates_6_ARLOCK;
  output [2:0] m_axi_updates_6_ARPROT;
  output [3:0] m_axi_updates_6_ARQOS;
  input m_axi_updates_6_ARREADY;
  output [3:0] m_axi_updates_6_ARREGION;
  output [2:0] m_axi_updates_6_ARSIZE;
  output m_axi_updates_6_ARUSER;
  output m_axi_updates_6_ARVALID;
  output [63:0] m_axi_updates_6_AWADDR;
  output [1:0] m_axi_updates_6_AWBURST;
  output [3:0] m_axi_updates_6_AWCACHE;
  output [0:0] m_axi_updates_6_AWID;
  output [7:0] m_axi_updates_6_AWLEN;
  output m_axi_updates_6_AWLOCK;
  output [2:0] m_axi_updates_6_AWPROT;
  output [3:0] m_axi_updates_6_AWQOS;
  input m_axi_updates_6_AWREADY;
  output [3:0] m_axi_updates_6_AWREGION;
  output [2:0] m_axi_updates_6_AWSIZE;
  output m_axi_updates_6_AWUSER;
  output m_axi_updates_6_AWVALID;
  input [0:0] m_axi_updates_6_BID;
  output m_axi_updates_6_BREADY;
  input [1:0] m_axi_updates_6_BRESP;
  input m_axi_updates_6_BUSER;
  input m_axi_updates_6_BVALID;
  input [511:0] m_axi_updates_6_RDATA;
  input [0:0] m_axi_updates_6_RID;
  input m_axi_updates_6_RLAST;
  output m_axi_updates_6_RREADY;
  input [1:0] m_axi_updates_6_RRESP;
  input m_axi_updates_6_RUSER;
  input m_axi_updates_6_RVALID;
  output [511:0] m_axi_updates_6_WDATA;
  output [0:0] m_axi_updates_6_WID;
  output m_axi_updates_6_WLAST;
  input m_axi_updates_6_WREADY;
  output [63:0] m_axi_updates_6_WSTRB;
  output m_axi_updates_6_WUSER;
  output m_axi_updates_6_WVALID;
  output [63:0] m_axi_updates_7_ARADDR;
  output [1:0] m_axi_updates_7_ARBURST;
  output [3:0] m_axi_updates_7_ARCACHE;
  output [0:0] m_axi_updates_7_ARID;
  output [7:0] m_axi_updates_7_ARLEN;
  output m_axi_updates_7_ARLOCK;
  output [2:0] m_axi_updates_7_ARPROT;
  output [3:0] m_axi_updates_7_ARQOS;
  input m_axi_updates_7_ARREADY;
  output [3:0] m_axi_updates_7_ARREGION;
  output [2:0] m_axi_updates_7_ARSIZE;
  output m_axi_updates_7_ARUSER;
  output m_axi_updates_7_ARVALID;
  output [63:0] m_axi_updates_7_AWADDR;
  output [1:0] m_axi_updates_7_AWBURST;
  output [3:0] m_axi_updates_7_AWCACHE;
  output [0:0] m_axi_updates_7_AWID;
  output [7:0] m_axi_updates_7_AWLEN;
  output m_axi_updates_7_AWLOCK;
  output [2:0] m_axi_updates_7_AWPROT;
  output [3:0] m_axi_updates_7_AWQOS;
  input m_axi_updates_7_AWREADY;
  output [3:0] m_axi_updates_7_AWREGION;
  output [2:0] m_axi_updates_7_AWSIZE;
  output m_axi_updates_7_AWUSER;
  output m_axi_updates_7_AWVALID;
  input [0:0] m_axi_updates_7_BID;
  output m_axi_updates_7_BREADY;
  input [1:0] m_axi_updates_7_BRESP;
  input m_axi_updates_7_BUSER;
  input m_axi_updates_7_BVALID;
  input [511:0] m_axi_updates_7_RDATA;
  input [0:0] m_axi_updates_7_RID;
  input m_axi_updates_7_RLAST;
  output m_axi_updates_7_RREADY;
  input [1:0] m_axi_updates_7_RRESP;
  input m_axi_updates_7_RUSER;
  input m_axi_updates_7_RVALID;
  output [511:0] m_axi_updates_7_WDATA;
  output [0:0] m_axi_updates_7_WID;
  output m_axi_updates_7_WLAST;
  input m_axi_updates_7_WREADY;
  output [63:0] m_axi_updates_7_WSTRB;
  output m_axi_updates_7_WUSER;
  output m_axi_updates_7_WVALID;
  output [63:0] m_axi_degrees_ARADDR;
  output [1:0] m_axi_degrees_ARBURST;
  output [3:0] m_axi_degrees_ARCACHE;
  output [0:0] m_axi_degrees_ARID;
  output [7:0] m_axi_degrees_ARLEN;
  output m_axi_degrees_ARLOCK;
  output [2:0] m_axi_degrees_ARPROT;
  output [3:0] m_axi_degrees_ARQOS;
  input m_axi_degrees_ARREADY;
  output [3:0] m_axi_degrees_ARREGION;
  output [2:0] m_axi_degrees_ARSIZE;
  output m_axi_degrees_ARUSER;
  output m_axi_degrees_ARVALID;
  output [63:0] m_axi_degrees_AWADDR;
  output [1:0] m_axi_degrees_AWBURST;
  output [3:0] m_axi_degrees_AWCACHE;
  output [0:0] m_axi_degrees_AWID;
  output [7:0] m_axi_degrees_AWLEN;
  output m_axi_degrees_AWLOCK;
  output [2:0] m_axi_degrees_AWPROT;
  output [3:0] m_axi_degrees_AWQOS;
  input m_axi_degrees_AWREADY;
  output [3:0] m_axi_degrees_AWREGION;
  output [2:0] m_axi_degrees_AWSIZE;
  output m_axi_degrees_AWUSER;
  output m_axi_degrees_AWVALID;
  input [0:0] m_axi_degrees_BID;
  output m_axi_degrees_BREADY;
  input [1:0] m_axi_degrees_BRESP;
  input m_axi_degrees_BUSER;
  input m_axi_degrees_BVALID;
  input [511:0] m_axi_degrees_RDATA;
  input [0:0] m_axi_degrees_RID;
  input m_axi_degrees_RLAST;
  output m_axi_degrees_RREADY;
  input [1:0] m_axi_degrees_RRESP;
  input m_axi_degrees_RUSER;
  input m_axi_degrees_RVALID;
  output [511:0] m_axi_degrees_WDATA;
  output [0:0] m_axi_degrees_WID;
  output m_axi_degrees_WLAST;
  input m_axi_degrees_WREADY;
  output [63:0] m_axi_degrees_WSTRB;
  output m_axi_degrees_WUSER;
  output m_axi_degrees_WVALID;
  output [63:0] m_axi_rankings_ARADDR;
  output [1:0] m_axi_rankings_ARBURST;
  output [3:0] m_axi_rankings_ARCACHE;
  output [0:0] m_axi_rankings_ARID;
  output [7:0] m_axi_rankings_ARLEN;
  output m_axi_rankings_ARLOCK;
  output [2:0] m_axi_rankings_ARPROT;
  output [3:0] m_axi_rankings_ARQOS;
  input m_axi_rankings_ARREADY;
  output [3:0] m_axi_rankings_ARREGION;
  output [2:0] m_axi_rankings_ARSIZE;
  output m_axi_rankings_ARUSER;
  output m_axi_rankings_ARVALID;
  output [63:0] m_axi_rankings_AWADDR;
  output [1:0] m_axi_rankings_AWBURST;
  output [3:0] m_axi_rankings_AWCACHE;
  output [0:0] m_axi_rankings_AWID;
  output [7:0] m_axi_rankings_AWLEN;
  output m_axi_rankings_AWLOCK;
  output [2:0] m_axi_rankings_AWPROT;
  output [3:0] m_axi_rankings_AWQOS;
  input m_axi_rankings_AWREADY;
  output [3:0] m_axi_rankings_AWREGION;
  output [2:0] m_axi_rankings_AWSIZE;
  output m_axi_rankings_AWUSER;
  output m_axi_rankings_AWVALID;
  input [0:0] m_axi_rankings_BID;
  output m_axi_rankings_BREADY;
  input [1:0] m_axi_rankings_BRESP;
  input m_axi_rankings_BUSER;
  input m_axi_rankings_BVALID;
  input [511:0] m_axi_rankings_RDATA;
  input [0:0] m_axi_rankings_RID;
  input m_axi_rankings_RLAST;
  output m_axi_rankings_RREADY;
  input [1:0] m_axi_rankings_RRESP;
  input m_axi_rankings_RUSER;
  input m_axi_rankings_RVALID;
  output [511:0] m_axi_rankings_WDATA;
  output [0:0] m_axi_rankings_WID;
  output m_axi_rankings_WLAST;
  input m_axi_rankings_WREADY;
  output [63:0] m_axi_rankings_WSTRB;
  output m_axi_rankings_WUSER;
  output m_axi_rankings_WVALID;
  output [63:0] m_axi_tmps_ARADDR;
  output [1:0] m_axi_tmps_ARBURST;
  output [3:0] m_axi_tmps_ARCACHE;
  output [0:0] m_axi_tmps_ARID;
  output [7:0] m_axi_tmps_ARLEN;
  output m_axi_tmps_ARLOCK;
  output [2:0] m_axi_tmps_ARPROT;
  output [3:0] m_axi_tmps_ARQOS;
  input m_axi_tmps_ARREADY;
  output [3:0] m_axi_tmps_ARREGION;
  output [2:0] m_axi_tmps_ARSIZE;
  output m_axi_tmps_ARUSER;
  output m_axi_tmps_ARVALID;
  output [63:0] m_axi_tmps_AWADDR;
  output [1:0] m_axi_tmps_AWBURST;
  output [3:0] m_axi_tmps_AWCACHE;
  output [0:0] m_axi_tmps_AWID;
  output [7:0] m_axi_tmps_AWLEN;
  output m_axi_tmps_AWLOCK;
  output [2:0] m_axi_tmps_AWPROT;
  output [3:0] m_axi_tmps_AWQOS;
  input m_axi_tmps_AWREADY;
  output [3:0] m_axi_tmps_AWREGION;
  output [2:0] m_axi_tmps_AWSIZE;
  output m_axi_tmps_AWUSER;
  output m_axi_tmps_AWVALID;
  input [0:0] m_axi_tmps_BID;
  output m_axi_tmps_BREADY;
  input [1:0] m_axi_tmps_BRESP;
  input m_axi_tmps_BUSER;
  input m_axi_tmps_BVALID;
  input [511:0] m_axi_tmps_RDATA;
  input [0:0] m_axi_tmps_RID;
  input m_axi_tmps_RLAST;
  output m_axi_tmps_RREADY;
  input [1:0] m_axi_tmps_RRESP;
  input m_axi_tmps_RUSER;
  input m_axi_tmps_RVALID;
  output [511:0] m_axi_tmps_WDATA;
  output [0:0] m_axi_tmps_WID;
  output m_axi_tmps_WLAST;
  input m_axi_tmps_WREADY;
  output [63:0] m_axi_tmps_WSTRB;
  output m_axi_tmps_WUSER;
  output m_axi_tmps_WVALID;
  wire ap_start;
  wire [15:0] num_partitions;
  wire [63:0] metadata;
  wire [63:0] degrees;
  wire [63:0] rankings;
  wire [63:0] tmps;
  wire [63:0] edges_0;
  wire [63:0] edges_1;
  wire [63:0] edges_2;
  wire [63:0] edges_3;
  wire [63:0] edges_4;
  wire [63:0] edges_5;
  wire [63:0] edges_6;
  wire [63:0] edges_7;
  wire [63:0] updates_0;
  wire [63:0] updates_1;
  wire [63:0] updates_2;
  wire [63:0] updates_3;
  wire [63:0] updates_4;
  wire [63:0] updates_5;
  wire [63:0] updates_6;
  wire [63:0] updates_7;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;
  wire ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg ap_rst_n__q2;
  wire [32:0] edge_req_0__dout;
  wire edge_req_0__empty_n;
  wire edge_req_0__read;
  wire [32:0] edge_req_0__din;
  wire edge_req_0__full_n;
  wire edge_req_0__write;
  wire edge_req_0__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_req_0__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_req_0__rst__q2;
  wire [32:0] edge_req_1__dout;
  wire edge_req_1__empty_n;
  wire edge_req_1__read;
  wire [32:0] edge_req_1__din;
  wire edge_req_1__full_n;
  wire edge_req_1__write;
  wire edge_req_1__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_req_1__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_req_1__rst__q2;
  wire [32:0] edge_req_2__dout;
  wire edge_req_2__empty_n;
  wire edge_req_2__read;
  wire [32:0] edge_req_2__din;
  wire edge_req_2__full_n;
  wire edge_req_2__write;
  wire edge_req_2__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_req_2__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_req_2__rst__q2;
  wire [32:0] edge_req_3__dout;
  wire edge_req_3__empty_n;
  wire edge_req_3__read;
  wire [32:0] edge_req_3__din;
  wire edge_req_3__full_n;
  wire edge_req_3__write;
  wire edge_req_3__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_req_3__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_req_3__rst__q2;
  wire [32:0] edge_req_4__dout;
  wire edge_req_4__empty_n;
  wire edge_req_4__read;
  wire [32:0] edge_req_4__din;
  wire edge_req_4__full_n;
  wire edge_req_4__write;
  wire edge_req_4__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_req_4__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_req_4__rst__q2;
  wire [32:0] edge_req_5__dout;
  wire edge_req_5__empty_n;
  wire edge_req_5__read;
  wire [32:0] edge_req_5__din;
  wire edge_req_5__full_n;
  wire edge_req_5__write;
  wire edge_req_5__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_req_5__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_req_5__rst__q2;
  wire [32:0] edge_req_6__dout;
  wire edge_req_6__empty_n;
  wire edge_req_6__read;
  wire [32:0] edge_req_6__din;
  wire edge_req_6__full_n;
  wire edge_req_6__write;
  wire edge_req_6__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_req_6__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_req_6__rst__q2;
  wire [32:0] edge_req_7__dout;
  wire edge_req_7__empty_n;
  wire edge_req_7__read;
  wire [32:0] edge_req_7__din;
  wire edge_req_7__full_n;
  wire edge_req_7__write;
  wire edge_req_7__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_req_7__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_req_7__rst__q2;
  wire [512:0] edge_resp_0__dout;
  wire edge_resp_0__empty_n;
  wire edge_resp_0__read;
  wire [512:0] edge_resp_0__din;
  wire edge_resp_0__full_n;
  wire edge_resp_0__write;
  wire edge_resp_0__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_resp_0__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_resp_0__rst__q2;
  wire [512:0] edge_resp_1__dout;
  wire edge_resp_1__empty_n;
  wire edge_resp_1__read;
  wire [512:0] edge_resp_1__din;
  wire edge_resp_1__full_n;
  wire edge_resp_1__write;
  wire edge_resp_1__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_resp_1__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_resp_1__rst__q2;
  wire [512:0] edge_resp_2__dout;
  wire edge_resp_2__empty_n;
  wire edge_resp_2__read;
  wire [512:0] edge_resp_2__din;
  wire edge_resp_2__full_n;
  wire edge_resp_2__write;
  wire edge_resp_2__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_resp_2__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_resp_2__rst__q2;
  wire [512:0] edge_resp_3__dout;
  wire edge_resp_3__empty_n;
  wire edge_resp_3__read;
  wire [512:0] edge_resp_3__din;
  wire edge_resp_3__full_n;
  wire edge_resp_3__write;
  wire edge_resp_3__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_resp_3__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_resp_3__rst__q2;
  wire [512:0] edge_resp_4__dout;
  wire edge_resp_4__empty_n;
  wire edge_resp_4__read;
  wire [512:0] edge_resp_4__din;
  wire edge_resp_4__full_n;
  wire edge_resp_4__write;
  wire edge_resp_4__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_resp_4__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_resp_4__rst__q2;
  wire [512:0] edge_resp_5__dout;
  wire edge_resp_5__empty_n;
  wire edge_resp_5__read;
  wire [512:0] edge_resp_5__din;
  wire edge_resp_5__full_n;
  wire edge_resp_5__write;
  wire edge_resp_5__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_resp_5__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_resp_5__rst__q2;
  wire [512:0] edge_resp_6__dout;
  wire edge_resp_6__empty_n;
  wire edge_resp_6__read;
  wire [512:0] edge_resp_6__din;
  wire edge_resp_6__full_n;
  wire edge_resp_6__write;
  wire edge_resp_6__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_resp_6__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_resp_6__rst__q2;
  wire [512:0] edge_resp_7__dout;
  wire edge_resp_7__empty_n;
  wire edge_resp_7__read;
  wire [512:0] edge_resp_7__din;
  wire edge_resp_7__full_n;
  wire edge_resp_7__write;
  wire edge_resp_7__rst__q0;
  (* dont_touch = "yes" *)
  reg edge_resp_7__rst__q1;
  (* dont_touch = "yes" *)
  reg edge_resp_7__rst__q2;
  wire [48:0] num_updates_0__dout;
  wire num_updates_0__empty_n;
  wire num_updates_0__read;
  wire [48:0] num_updates_0__din;
  wire num_updates_0__full_n;
  wire num_updates_0__write;
  wire num_updates_0__rst__q0;
  (* dont_touch = "yes" *)
  reg num_updates_0__rst__q1;
  (* dont_touch = "yes" *)
  reg num_updates_0__rst__q2;
  wire [48:0] num_updates_1__dout;
  wire num_updates_1__empty_n;
  wire num_updates_1__read;
  wire [48:0] num_updates_1__din;
  wire num_updates_1__full_n;
  wire num_updates_1__write;
  wire num_updates_1__rst__q0;
  (* dont_touch = "yes" *)
  reg num_updates_1__rst__q1;
  (* dont_touch = "yes" *)
  reg num_updates_1__rst__q2;
  wire [48:0] num_updates_2__dout;
  wire num_updates_2__empty_n;
  wire num_updates_2__read;
  wire [48:0] num_updates_2__din;
  wire num_updates_2__full_n;
  wire num_updates_2__write;
  wire num_updates_2__rst__q0;
  (* dont_touch = "yes" *)
  reg num_updates_2__rst__q1;
  (* dont_touch = "yes" *)
  reg num_updates_2__rst__q2;
  wire [48:0] num_updates_3__dout;
  wire num_updates_3__empty_n;
  wire num_updates_3__read;
  wire [48:0] num_updates_3__din;
  wire num_updates_3__full_n;
  wire num_updates_3__write;
  wire num_updates_3__rst__q0;
  (* dont_touch = "yes" *)
  reg num_updates_3__rst__q1;
  (* dont_touch = "yes" *)
  reg num_updates_3__rst__q2;
  wire [48:0] num_updates_4__dout;
  wire num_updates_4__empty_n;
  wire num_updates_4__read;
  wire [48:0] num_updates_4__din;
  wire num_updates_4__full_n;
  wire num_updates_4__write;
  wire num_updates_4__rst__q0;
  (* dont_touch = "yes" *)
  reg num_updates_4__rst__q1;
  (* dont_touch = "yes" *)
  reg num_updates_4__rst__q2;
  wire [48:0] num_updates_5__dout;
  wire num_updates_5__empty_n;
  wire num_updates_5__read;
  wire [48:0] num_updates_5__din;
  wire num_updates_5__full_n;
  wire num_updates_5__write;
  wire num_updates_5__rst__q0;
  (* dont_touch = "yes" *)
  reg num_updates_5__rst__q1;
  (* dont_touch = "yes" *)
  reg num_updates_5__rst__q2;
  wire [48:0] num_updates_6__dout;
  wire num_updates_6__empty_n;
  wire num_updates_6__read;
  wire [48:0] num_updates_6__din;
  wire num_updates_6__full_n;
  wire num_updates_6__write;
  wire num_updates_6__rst__q0;
  (* dont_touch = "yes" *)
  reg num_updates_6__rst__q1;
  (* dont_touch = "yes" *)
  reg num_updates_6__rst__q2;
  wire [48:0] num_updates_7__dout;
  wire num_updates_7__empty_n;
  wire num_updates_7__read;
  wire [48:0] num_updates_7__din;
  wire num_updates_7__full_n;
  wire num_updates_7__write;
  wire num_updates_7__rst__q0;
  (* dont_touch = "yes" *)
  reg num_updates_7__rst__q1;
  (* dont_touch = "yes" *)
  reg num_updates_7__rst__q2;
  wire [64:0] scatter_phase_vertex_req__dout;
  wire scatter_phase_vertex_req__empty_n;
  wire scatter_phase_vertex_req__read;
  wire [64:0] scatter_phase_vertex_req__din;
  wire scatter_phase_vertex_req__full_n;
  wire scatter_phase_vertex_req__write;
  wire scatter_phase_vertex_req__rst__q0;
  (* dont_touch = "yes" *)
  reg scatter_phase_vertex_req__rst__q1;
  (* dont_touch = "yes" *)
  reg scatter_phase_vertex_req__rst__q2;
  wire [210:0] task_req_0__dout;
  wire task_req_0__empty_n;
  wire task_req_0__read;
  wire [210:0] task_req_0__din;
  wire task_req_0__full_n;
  wire task_req_0__write;
  wire task_req_0__rst__q0;
  (* dont_touch = "yes" *)
  reg task_req_0__rst__q1;
  (* dont_touch = "yes" *)
  reg task_req_0__rst__q2;
  wire [210:0] task_req_1__dout;
  wire task_req_1__empty_n;
  wire task_req_1__read;
  wire [210:0] task_req_1__din;
  wire task_req_1__full_n;
  wire task_req_1__write;
  wire task_req_1__rst__q0;
  (* dont_touch = "yes" *)
  reg task_req_1__rst__q1;
  (* dont_touch = "yes" *)
  reg task_req_1__rst__q2;
  wire [210:0] task_req_2__dout;
  wire task_req_2__empty_n;
  wire task_req_2__read;
  wire [210:0] task_req_2__din;
  wire task_req_2__full_n;
  wire task_req_2__write;
  wire task_req_2__rst__q0;
  (* dont_touch = "yes" *)
  reg task_req_2__rst__q1;
  (* dont_touch = "yes" *)
  reg task_req_2__rst__q2;
  wire [210:0] task_req_3__dout;
  wire task_req_3__empty_n;
  wire task_req_3__read;
  wire [210:0] task_req_3__din;
  wire task_req_3__full_n;
  wire task_req_3__write;
  wire task_req_3__rst__q0;
  (* dont_touch = "yes" *)
  reg task_req_3__rst__q1;
  (* dont_touch = "yes" *)
  reg task_req_3__rst__q2;
  wire [210:0] task_req_4__dout;
  wire task_req_4__empty_n;
  wire task_req_4__read;
  wire [210:0] task_req_4__din;
  wire task_req_4__full_n;
  wire task_req_4__write;
  wire task_req_4__rst__q0;
  (* dont_touch = "yes" *)
  reg task_req_4__rst__q1;
  (* dont_touch = "yes" *)
  reg task_req_4__rst__q2;
  wire [210:0] task_req_5__dout;
  wire task_req_5__empty_n;
  wire task_req_5__read;
  wire [210:0] task_req_5__din;
  wire task_req_5__full_n;
  wire task_req_5__write;
  wire task_req_5__rst__q0;
  (* dont_touch = "yes" *)
  reg task_req_5__rst__q1;
  (* dont_touch = "yes" *)
  reg task_req_5__rst__q2;
  wire [210:0] task_req_6__dout;
  wire task_req_6__empty_n;
  wire task_req_6__read;
  wire [210:0] task_req_6__din;
  wire task_req_6__full_n;
  wire task_req_6__write;
  wire task_req_6__rst__q0;
  (* dont_touch = "yes" *)
  reg task_req_6__rst__q1;
  (* dont_touch = "yes" *)
  reg task_req_6__rst__q2;
  wire [210:0] task_req_7__dout;
  wire task_req_7__empty_n;
  wire task_req_7__read;
  wire [210:0] task_req_7__din;
  wire task_req_7__full_n;
  wire task_req_7__write;
  wire task_req_7__rst__q0;
  (* dont_touch = "yes" *)
  reg task_req_7__rst__q1;
  (* dont_touch = "yes" *)
  reg task_req_7__rst__q2;
  wire [1:0] task_resp_0__dout;
  wire task_resp_0__empty_n;
  wire task_resp_0__read;
  wire [1:0] task_resp_0__din;
  wire task_resp_0__full_n;
  wire task_resp_0__write;
  wire task_resp_0__rst__q0;
  (* dont_touch = "yes" *)
  reg task_resp_0__rst__q1;
  (* dont_touch = "yes" *)
  reg task_resp_0__rst__q2;
  wire [1:0] task_resp_1__dout;
  wire task_resp_1__empty_n;
  wire task_resp_1__read;
  wire [1:0] task_resp_1__din;
  wire task_resp_1__full_n;
  wire task_resp_1__write;
  wire task_resp_1__rst__q0;
  (* dont_touch = "yes" *)
  reg task_resp_1__rst__q1;
  (* dont_touch = "yes" *)
  reg task_resp_1__rst__q2;
  wire [1:0] task_resp_2__dout;
  wire task_resp_2__empty_n;
  wire task_resp_2__read;
  wire [1:0] task_resp_2__din;
  wire task_resp_2__full_n;
  wire task_resp_2__write;
  wire task_resp_2__rst__q0;
  (* dont_touch = "yes" *)
  reg task_resp_2__rst__q1;
  (* dont_touch = "yes" *)
  reg task_resp_2__rst__q2;
  wire [1:0] task_resp_3__dout;
  wire task_resp_3__empty_n;
  wire task_resp_3__read;
  wire [1:0] task_resp_3__din;
  wire task_resp_3__full_n;
  wire task_resp_3__write;
  wire task_resp_3__rst__q0;
  (* dont_touch = "yes" *)
  reg task_resp_3__rst__q1;
  (* dont_touch = "yes" *)
  reg task_resp_3__rst__q2;
  wire [1:0] task_resp_4__dout;
  wire task_resp_4__empty_n;
  wire task_resp_4__read;
  wire [1:0] task_resp_4__din;
  wire task_resp_4__full_n;
  wire task_resp_4__write;
  wire task_resp_4__rst__q0;
  (* dont_touch = "yes" *)
  reg task_resp_4__rst__q1;
  (* dont_touch = "yes" *)
  reg task_resp_4__rst__q2;
  wire [1:0] task_resp_5__dout;
  wire task_resp_5__empty_n;
  wire task_resp_5__read;
  wire [1:0] task_resp_5__din;
  wire task_resp_5__full_n;
  wire task_resp_5__write;
  wire task_resp_5__rst__q0;
  (* dont_touch = "yes" *)
  reg task_resp_5__rst__q1;
  (* dont_touch = "yes" *)
  reg task_resp_5__rst__q2;
  wire [1:0] task_resp_6__dout;
  wire task_resp_6__empty_n;
  wire task_resp_6__read;
  wire [1:0] task_resp_6__din;
  wire task_resp_6__full_n;
  wire task_resp_6__write;
  wire task_resp_6__rst__q0;
  (* dont_touch = "yes" *)
  reg task_resp_6__rst__q1;
  (* dont_touch = "yes" *)
  reg task_resp_6__rst__q2;
  wire [1:0] task_resp_7__dout;
  wire task_resp_7__empty_n;
  wire task_resp_7__read;
  wire [1:0] task_resp_7__din;
  wire task_resp_7__full_n;
  wire task_resp_7__write;
  wire task_resp_7__rst__q0;
  (* dont_touch = "yes" *)
  reg task_resp_7__rst__q1;
  (* dont_touch = "yes" *)
  reg task_resp_7__rst__q2;
  wire [32:0] update_config_0__dout;
  wire update_config_0__empty_n;
  wire update_config_0__read;
  wire [32:0] update_config_0__din;
  wire update_config_0__full_n;
  wire update_config_0__write;
  wire update_config_0__rst__q0;
  (* dont_touch = "yes" *)
  reg update_config_0__rst__q1;
  (* dont_touch = "yes" *)
  reg update_config_0__rst__q2;
  wire [32:0] update_config_1__dout;
  wire update_config_1__empty_n;
  wire update_config_1__read;
  wire [32:0] update_config_1__din;
  wire update_config_1__full_n;
  wire update_config_1__write;
  wire update_config_1__rst__q0;
  (* dont_touch = "yes" *)
  reg update_config_1__rst__q1;
  (* dont_touch = "yes" *)
  reg update_config_1__rst__q2;
  wire [32:0] update_config_2__dout;
  wire update_config_2__empty_n;
  wire update_config_2__read;
  wire [32:0] update_config_2__din;
  wire update_config_2__full_n;
  wire update_config_2__write;
  wire update_config_2__rst__q0;
  (* dont_touch = "yes" *)
  reg update_config_2__rst__q1;
  (* dont_touch = "yes" *)
  reg update_config_2__rst__q2;
  wire [32:0] update_config_3__dout;
  wire update_config_3__empty_n;
  wire update_config_3__read;
  wire [32:0] update_config_3__din;
  wire update_config_3__full_n;
  wire update_config_3__write;
  wire update_config_3__rst__q0;
  (* dont_touch = "yes" *)
  reg update_config_3__rst__q1;
  (* dont_touch = "yes" *)
  reg update_config_3__rst__q2;
  wire [32:0] update_config_4__dout;
  wire update_config_4__empty_n;
  wire update_config_4__read;
  wire [32:0] update_config_4__din;
  wire update_config_4__full_n;
  wire update_config_4__write;
  wire update_config_4__rst__q0;
  (* dont_touch = "yes" *)
  reg update_config_4__rst__q1;
  (* dont_touch = "yes" *)
  reg update_config_4__rst__q2;
  wire [32:0] update_config_5__dout;
  wire update_config_5__empty_n;
  wire update_config_5__read;
  wire [32:0] update_config_5__din;
  wire update_config_5__full_n;
  wire update_config_5__write;
  wire update_config_5__rst__q0;
  (* dont_touch = "yes" *)
  reg update_config_5__rst__q1;
  (* dont_touch = "yes" *)
  reg update_config_5__rst__q2;
  wire [32:0] update_config_6__dout;
  wire update_config_6__empty_n;
  wire update_config_6__read;
  wire [32:0] update_config_6__din;
  wire update_config_6__full_n;
  wire update_config_6__write;
  wire update_config_6__rst__q0;
  (* dont_touch = "yes" *)
  reg update_config_6__rst__q1;
  (* dont_touch = "yes" *)
  reg update_config_6__rst__q2;
  wire [32:0] update_config_7__dout;
  wire update_config_7__empty_n;
  wire update_config_7__read;
  wire [32:0] update_config_7__din;
  wire update_config_7__full_n;
  wire update_config_7__write;
  wire update_config_7__rst__q0;
  (* dont_touch = "yes" *)
  reg update_config_7__rst__q1;
  (* dont_touch = "yes" *)
  reg update_config_7__rst__q2;
  wire [512:0] update_mm2pe_0__dout;
  wire update_mm2pe_0__empty_n;
  wire update_mm2pe_0__read;
  wire [512:0] update_mm2pe_0__din;
  wire update_mm2pe_0__full_n;
  wire update_mm2pe_0__write;
  wire update_mm2pe_0__rst__q0;
  (* dont_touch = "yes" *)
  reg update_mm2pe_0__rst__q1;
  (* dont_touch = "yes" *)
  reg update_mm2pe_0__rst__q2;
  wire [512:0] update_mm2pe_1__dout;
  wire update_mm2pe_1__empty_n;
  wire update_mm2pe_1__read;
  wire [512:0] update_mm2pe_1__din;
  wire update_mm2pe_1__full_n;
  wire update_mm2pe_1__write;
  wire update_mm2pe_1__rst__q0;
  (* dont_touch = "yes" *)
  reg update_mm2pe_1__rst__q1;
  (* dont_touch = "yes" *)
  reg update_mm2pe_1__rst__q2;
  wire [512:0] update_mm2pe_2__dout;
  wire update_mm2pe_2__empty_n;
  wire update_mm2pe_2__read;
  wire [512:0] update_mm2pe_2__din;
  wire update_mm2pe_2__full_n;
  wire update_mm2pe_2__write;
  wire update_mm2pe_2__rst__q0;
  (* dont_touch = "yes" *)
  reg update_mm2pe_2__rst__q1;
  (* dont_touch = "yes" *)
  reg update_mm2pe_2__rst__q2;
  wire [512:0] update_mm2pe_3__dout;
  wire update_mm2pe_3__empty_n;
  wire update_mm2pe_3__read;
  wire [512:0] update_mm2pe_3__din;
  wire update_mm2pe_3__full_n;
  wire update_mm2pe_3__write;
  wire update_mm2pe_3__rst__q0;
  (* dont_touch = "yes" *)
  reg update_mm2pe_3__rst__q1;
  (* dont_touch = "yes" *)
  reg update_mm2pe_3__rst__q2;
  wire [512:0] update_mm2pe_4__dout;
  wire update_mm2pe_4__empty_n;
  wire update_mm2pe_4__read;
  wire [512:0] update_mm2pe_4__din;
  wire update_mm2pe_4__full_n;
  wire update_mm2pe_4__write;
  wire update_mm2pe_4__rst__q0;
  (* dont_touch = "yes" *)
  reg update_mm2pe_4__rst__q1;
  (* dont_touch = "yes" *)
  reg update_mm2pe_4__rst__q2;
  wire [512:0] update_mm2pe_5__dout;
  wire update_mm2pe_5__empty_n;
  wire update_mm2pe_5__read;
  wire [512:0] update_mm2pe_5__din;
  wire update_mm2pe_5__full_n;
  wire update_mm2pe_5__write;
  wire update_mm2pe_5__rst__q0;
  (* dont_touch = "yes" *)
  reg update_mm2pe_5__rst__q1;
  (* dont_touch = "yes" *)
  reg update_mm2pe_5__rst__q2;
  wire [512:0] update_mm2pe_6__dout;
  wire update_mm2pe_6__empty_n;
  wire update_mm2pe_6__read;
  wire [512:0] update_mm2pe_6__din;
  wire update_mm2pe_6__full_n;
  wire update_mm2pe_6__write;
  wire update_mm2pe_6__rst__q0;
  (* dont_touch = "yes" *)
  reg update_mm2pe_6__rst__q1;
  (* dont_touch = "yes" *)
  reg update_mm2pe_6__rst__q2;
  wire [512:0] update_mm2pe_7__dout;
  wire update_mm2pe_7__empty_n;
  wire update_mm2pe_7__read;
  wire [512:0] update_mm2pe_7__din;
  wire update_mm2pe_7__full_n;
  wire update_mm2pe_7__write;
  wire update_mm2pe_7__rst__q0;
  (* dont_touch = "yes" *)
  reg update_mm2pe_7__rst__q1;
  (* dont_touch = "yes" *)
  reg update_mm2pe_7__rst__q2;
  wire [528:0] update_pe2mm_0__dout;
  wire update_pe2mm_0__empty_n;
  wire update_pe2mm_0__read;
  wire [528:0] update_pe2mm_0__din;
  wire update_pe2mm_0__full_n;
  wire update_pe2mm_0__write;
  wire update_pe2mm_0__rst__q0;
  (* dont_touch = "yes" *)
  reg update_pe2mm_0__rst__q1;
  (* dont_touch = "yes" *)
  reg update_pe2mm_0__rst__q2;
  wire [528:0] update_pe2mm_1__dout;
  wire update_pe2mm_1__empty_n;
  wire update_pe2mm_1__read;
  wire [528:0] update_pe2mm_1__din;
  wire update_pe2mm_1__full_n;
  wire update_pe2mm_1__write;
  wire update_pe2mm_1__rst__q0;
  (* dont_touch = "yes" *)
  reg update_pe2mm_1__rst__q1;
  (* dont_touch = "yes" *)
  reg update_pe2mm_1__rst__q2;
  wire [528:0] update_pe2mm_2__dout;
  wire update_pe2mm_2__empty_n;
  wire update_pe2mm_2__read;
  wire [528:0] update_pe2mm_2__din;
  wire update_pe2mm_2__full_n;
  wire update_pe2mm_2__write;
  wire update_pe2mm_2__rst__q0;
  (* dont_touch = "yes" *)
  reg update_pe2mm_2__rst__q1;
  (* dont_touch = "yes" *)
  reg update_pe2mm_2__rst__q2;
  wire [528:0] update_pe2mm_3__dout;
  wire update_pe2mm_3__empty_n;
  wire update_pe2mm_3__read;
  wire [528:0] update_pe2mm_3__din;
  wire update_pe2mm_3__full_n;
  wire update_pe2mm_3__write;
  wire update_pe2mm_3__rst__q0;
  (* dont_touch = "yes" *)
  reg update_pe2mm_3__rst__q1;
  (* dont_touch = "yes" *)
  reg update_pe2mm_3__rst__q2;
  wire [528:0] update_pe2mm_4__dout;
  wire update_pe2mm_4__empty_n;
  wire update_pe2mm_4__read;
  wire [528:0] update_pe2mm_4__din;
  wire update_pe2mm_4__full_n;
  wire update_pe2mm_4__write;
  wire update_pe2mm_4__rst__q0;
  (* dont_touch = "yes" *)
  reg update_pe2mm_4__rst__q1;
  (* dont_touch = "yes" *)
  reg update_pe2mm_4__rst__q2;
  wire [528:0] update_pe2mm_5__dout;
  wire update_pe2mm_5__empty_n;
  wire update_pe2mm_5__read;
  wire [528:0] update_pe2mm_5__din;
  wire update_pe2mm_5__full_n;
  wire update_pe2mm_5__write;
  wire update_pe2mm_5__rst__q0;
  (* dont_touch = "yes" *)
  reg update_pe2mm_5__rst__q1;
  (* dont_touch = "yes" *)
  reg update_pe2mm_5__rst__q2;
  wire [528:0] update_pe2mm_6__dout;
  wire update_pe2mm_6__empty_n;
  wire update_pe2mm_6__read;
  wire [528:0] update_pe2mm_6__din;
  wire update_pe2mm_6__full_n;
  wire update_pe2mm_6__write;
  wire update_pe2mm_6__rst__q0;
  (* dont_touch = "yes" *)
  reg update_pe2mm_6__rst__q1;
  (* dont_touch = "yes" *)
  reg update_pe2mm_6__rst__q2;
  wire [528:0] update_pe2mm_7__dout;
  wire update_pe2mm_7__empty_n;
  wire update_pe2mm_7__read;
  wire [528:0] update_pe2mm_7__din;
  wire update_pe2mm_7__full_n;
  wire update_pe2mm_7__write;
  wire update_pe2mm_7__rst__q0;
  (* dont_touch = "yes" *)
  reg update_pe2mm_7__rst__q1;
  (* dont_touch = "yes" *)
  reg update_pe2mm_7__rst__q2;
  wire [1:0] update_phase_0__dout;
  wire update_phase_0__empty_n;
  wire update_phase_0__read;
  wire [1:0] update_phase_0__din;
  wire update_phase_0__full_n;
  wire update_phase_0__write;
  wire update_phase_0__rst__q0;
  (* dont_touch = "yes" *)
  reg update_phase_0__rst__q1;
  (* dont_touch = "yes" *)
  reg update_phase_0__rst__q2;
  wire [1:0] update_phase_1__dout;
  wire update_phase_1__empty_n;
  wire update_phase_1__read;
  wire [1:0] update_phase_1__din;
  wire update_phase_1__full_n;
  wire update_phase_1__write;
  wire update_phase_1__rst__q0;
  (* dont_touch = "yes" *)
  reg update_phase_1__rst__q1;
  (* dont_touch = "yes" *)
  reg update_phase_1__rst__q2;
  wire [1:0] update_phase_2__dout;
  wire update_phase_2__empty_n;
  wire update_phase_2__read;
  wire [1:0] update_phase_2__din;
  wire update_phase_2__full_n;
  wire update_phase_2__write;
  wire update_phase_2__rst__q0;
  (* dont_touch = "yes" *)
  reg update_phase_2__rst__q1;
  (* dont_touch = "yes" *)
  reg update_phase_2__rst__q2;
  wire [1:0] update_phase_3__dout;
  wire update_phase_3__empty_n;
  wire update_phase_3__read;
  wire [1:0] update_phase_3__din;
  wire update_phase_3__full_n;
  wire update_phase_3__write;
  wire update_phase_3__rst__q0;
  (* dont_touch = "yes" *)
  reg update_phase_3__rst__q1;
  (* dont_touch = "yes" *)
  reg update_phase_3__rst__q2;
  wire [1:0] update_phase_4__dout;
  wire update_phase_4__empty_n;
  wire update_phase_4__read;
  wire [1:0] update_phase_4__din;
  wire update_phase_4__full_n;
  wire update_phase_4__write;
  wire update_phase_4__rst__q0;
  (* dont_touch = "yes" *)
  reg update_phase_4__rst__q1;
  (* dont_touch = "yes" *)
  reg update_phase_4__rst__q2;
  wire [1:0] update_phase_5__dout;
  wire update_phase_5__empty_n;
  wire update_phase_5__read;
  wire [1:0] update_phase_5__din;
  wire update_phase_5__full_n;
  wire update_phase_5__write;
  wire update_phase_5__rst__q0;
  (* dont_touch = "yes" *)
  reg update_phase_5__rst__q1;
  (* dont_touch = "yes" *)
  reg update_phase_5__rst__q2;
  wire [1:0] update_phase_6__dout;
  wire update_phase_6__empty_n;
  wire update_phase_6__read;
  wire [1:0] update_phase_6__din;
  wire update_phase_6__full_n;
  wire update_phase_6__write;
  wire update_phase_6__rst__q0;
  (* dont_touch = "yes" *)
  reg update_phase_6__rst__q1;
  (* dont_touch = "yes" *)
  reg update_phase_6__rst__q2;
  wire [1:0] update_phase_7__dout;
  wire update_phase_7__empty_n;
  wire update_phase_7__read;
  wire [1:0] update_phase_7__din;
  wire update_phase_7__full_n;
  wire update_phase_7__write;
  wire update_phase_7__rst__q0;
  (* dont_touch = "yes" *)
  reg update_phase_7__rst__q1;
  (* dont_touch = "yes" *)
  reg update_phase_7__rst__q2;
  wire [64:0] update_read_addr_0__dout;
  wire update_read_addr_0__empty_n;
  wire update_read_addr_0__read;
  wire [64:0] update_read_addr_0__din;
  wire update_read_addr_0__full_n;
  wire update_read_addr_0__write;
  wire update_read_addr_0__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_addr_0__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_addr_0__rst__q2;
  wire [64:0] update_read_addr_1__dout;
  wire update_read_addr_1__empty_n;
  wire update_read_addr_1__read;
  wire [64:0] update_read_addr_1__din;
  wire update_read_addr_1__full_n;
  wire update_read_addr_1__write;
  wire update_read_addr_1__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_addr_1__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_addr_1__rst__q2;
  wire [64:0] update_read_addr_2__dout;
  wire update_read_addr_2__empty_n;
  wire update_read_addr_2__read;
  wire [64:0] update_read_addr_2__din;
  wire update_read_addr_2__full_n;
  wire update_read_addr_2__write;
  wire update_read_addr_2__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_addr_2__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_addr_2__rst__q2;
  wire [64:0] update_read_addr_3__dout;
  wire update_read_addr_3__empty_n;
  wire update_read_addr_3__read;
  wire [64:0] update_read_addr_3__din;
  wire update_read_addr_3__full_n;
  wire update_read_addr_3__write;
  wire update_read_addr_3__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_addr_3__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_addr_3__rst__q2;
  wire [64:0] update_read_addr_4__dout;
  wire update_read_addr_4__empty_n;
  wire update_read_addr_4__read;
  wire [64:0] update_read_addr_4__din;
  wire update_read_addr_4__full_n;
  wire update_read_addr_4__write;
  wire update_read_addr_4__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_addr_4__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_addr_4__rst__q2;
  wire [64:0] update_read_addr_5__dout;
  wire update_read_addr_5__empty_n;
  wire update_read_addr_5__read;
  wire [64:0] update_read_addr_5__din;
  wire update_read_addr_5__full_n;
  wire update_read_addr_5__write;
  wire update_read_addr_5__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_addr_5__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_addr_5__rst__q2;
  wire [64:0] update_read_addr_6__dout;
  wire update_read_addr_6__empty_n;
  wire update_read_addr_6__read;
  wire [64:0] update_read_addr_6__din;
  wire update_read_addr_6__full_n;
  wire update_read_addr_6__write;
  wire update_read_addr_6__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_addr_6__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_addr_6__rst__q2;
  wire [64:0] update_read_addr_7__dout;
  wire update_read_addr_7__empty_n;
  wire update_read_addr_7__read;
  wire [64:0] update_read_addr_7__din;
  wire update_read_addr_7__full_n;
  wire update_read_addr_7__write;
  wire update_read_addr_7__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_addr_7__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_addr_7__rst__q2;
  wire [512:0] update_read_data_0__dout;
  wire update_read_data_0__empty_n;
  wire update_read_data_0__read;
  wire [512:0] update_read_data_0__din;
  wire update_read_data_0__full_n;
  wire update_read_data_0__write;
  wire update_read_data_0__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_data_0__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_data_0__rst__q2;
  wire [512:0] update_read_data_1__dout;
  wire update_read_data_1__empty_n;
  wire update_read_data_1__read;
  wire [512:0] update_read_data_1__din;
  wire update_read_data_1__full_n;
  wire update_read_data_1__write;
  wire update_read_data_1__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_data_1__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_data_1__rst__q2;
  wire [512:0] update_read_data_2__dout;
  wire update_read_data_2__empty_n;
  wire update_read_data_2__read;
  wire [512:0] update_read_data_2__din;
  wire update_read_data_2__full_n;
  wire update_read_data_2__write;
  wire update_read_data_2__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_data_2__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_data_2__rst__q2;
  wire [512:0] update_read_data_3__dout;
  wire update_read_data_3__empty_n;
  wire update_read_data_3__read;
  wire [512:0] update_read_data_3__din;
  wire update_read_data_3__full_n;
  wire update_read_data_3__write;
  wire update_read_data_3__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_data_3__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_data_3__rst__q2;
  wire [512:0] update_read_data_4__dout;
  wire update_read_data_4__empty_n;
  wire update_read_data_4__read;
  wire [512:0] update_read_data_4__din;
  wire update_read_data_4__full_n;
  wire update_read_data_4__write;
  wire update_read_data_4__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_data_4__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_data_4__rst__q2;
  wire [512:0] update_read_data_5__dout;
  wire update_read_data_5__empty_n;
  wire update_read_data_5__read;
  wire [512:0] update_read_data_5__din;
  wire update_read_data_5__full_n;
  wire update_read_data_5__write;
  wire update_read_data_5__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_data_5__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_data_5__rst__q2;
  wire [512:0] update_read_data_6__dout;
  wire update_read_data_6__empty_n;
  wire update_read_data_6__read;
  wire [512:0] update_read_data_6__din;
  wire update_read_data_6__full_n;
  wire update_read_data_6__write;
  wire update_read_data_6__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_data_6__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_data_6__rst__q2;
  wire [512:0] update_read_data_7__dout;
  wire update_read_data_7__empty_n;
  wire update_read_data_7__read;
  wire [512:0] update_read_data_7__din;
  wire update_read_data_7__full_n;
  wire update_read_data_7__write;
  wire update_read_data_7__rst__q0;
  (* dont_touch = "yes" *)
  reg update_read_data_7__rst__q1;
  (* dont_touch = "yes" *)
  reg update_read_data_7__rst__q2;
  wire [49:0] update_req_0__dout;
  wire update_req_0__empty_n;
  wire update_req_0__read;
  wire [49:0] update_req_0__din;
  wire update_req_0__full_n;
  wire update_req_0__write;
  wire update_req_0__rst__q0;
  (* dont_touch = "yes" *)
  reg update_req_0__rst__q1;
  (* dont_touch = "yes" *)
  reg update_req_0__rst__q2;
  wire [49:0] update_req_1__dout;
  wire update_req_1__empty_n;
  wire update_req_1__read;
  wire [49:0] update_req_1__din;
  wire update_req_1__full_n;
  wire update_req_1__write;
  wire update_req_1__rst__q0;
  (* dont_touch = "yes" *)
  reg update_req_1__rst__q1;
  (* dont_touch = "yes" *)
  reg update_req_1__rst__q2;
  wire [49:0] update_req_2__dout;
  wire update_req_2__empty_n;
  wire update_req_2__read;
  wire [49:0] update_req_2__din;
  wire update_req_2__full_n;
  wire update_req_2__write;
  wire update_req_2__rst__q0;
  (* dont_touch = "yes" *)
  reg update_req_2__rst__q1;
  (* dont_touch = "yes" *)
  reg update_req_2__rst__q2;
  wire [49:0] update_req_3__dout;
  wire update_req_3__empty_n;
  wire update_req_3__read;
  wire [49:0] update_req_3__din;
  wire update_req_3__full_n;
  wire update_req_3__write;
  wire update_req_3__rst__q0;
  (* dont_touch = "yes" *)
  reg update_req_3__rst__q1;
  (* dont_touch = "yes" *)
  reg update_req_3__rst__q2;
  wire [49:0] update_req_4__dout;
  wire update_req_4__empty_n;
  wire update_req_4__read;
  wire [49:0] update_req_4__din;
  wire update_req_4__full_n;
  wire update_req_4__write;
  wire update_req_4__rst__q0;
  (* dont_touch = "yes" *)
  reg update_req_4__rst__q1;
  (* dont_touch = "yes" *)
  reg update_req_4__rst__q2;
  wire [49:0] update_req_5__dout;
  wire update_req_5__empty_n;
  wire update_req_5__read;
  wire [49:0] update_req_5__din;
  wire update_req_5__full_n;
  wire update_req_5__write;
  wire update_req_5__rst__q0;
  (* dont_touch = "yes" *)
  reg update_req_5__rst__q1;
  (* dont_touch = "yes" *)
  reg update_req_5__rst__q2;
  wire [49:0] update_req_6__dout;
  wire update_req_6__empty_n;
  wire update_req_6__read;
  wire [49:0] update_req_6__din;
  wire update_req_6__full_n;
  wire update_req_6__write;
  wire update_req_6__rst__q0;
  (* dont_touch = "yes" *)
  reg update_req_6__rst__q1;
  (* dont_touch = "yes" *)
  reg update_req_6__rst__q2;
  wire [49:0] update_req_7__dout;
  wire update_req_7__empty_n;
  wire update_req_7__read;
  wire [49:0] update_req_7__din;
  wire update_req_7__full_n;
  wire update_req_7__write;
  wire update_req_7__rst__q0;
  (* dont_touch = "yes" *)
  reg update_req_7__rst__q1;
  (* dont_touch = "yes" *)
  reg update_req_7__rst__q2;
  wire [64:0] update_write_addr_0__dout;
  wire update_write_addr_0__empty_n;
  wire update_write_addr_0__read;
  wire [64:0] update_write_addr_0__din;
  wire update_write_addr_0__full_n;
  wire update_write_addr_0__write;
  wire update_write_addr_0__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_addr_0__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_addr_0__rst__q2;
  wire [64:0] update_write_addr_1__dout;
  wire update_write_addr_1__empty_n;
  wire update_write_addr_1__read;
  wire [64:0] update_write_addr_1__din;
  wire update_write_addr_1__full_n;
  wire update_write_addr_1__write;
  wire update_write_addr_1__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_addr_1__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_addr_1__rst__q2;
  wire [64:0] update_write_addr_2__dout;
  wire update_write_addr_2__empty_n;
  wire update_write_addr_2__read;
  wire [64:0] update_write_addr_2__din;
  wire update_write_addr_2__full_n;
  wire update_write_addr_2__write;
  wire update_write_addr_2__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_addr_2__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_addr_2__rst__q2;
  wire [64:0] update_write_addr_3__dout;
  wire update_write_addr_3__empty_n;
  wire update_write_addr_3__read;
  wire [64:0] update_write_addr_3__din;
  wire update_write_addr_3__full_n;
  wire update_write_addr_3__write;
  wire update_write_addr_3__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_addr_3__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_addr_3__rst__q2;
  wire [64:0] update_write_addr_4__dout;
  wire update_write_addr_4__empty_n;
  wire update_write_addr_4__read;
  wire [64:0] update_write_addr_4__din;
  wire update_write_addr_4__full_n;
  wire update_write_addr_4__write;
  wire update_write_addr_4__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_addr_4__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_addr_4__rst__q2;
  wire [64:0] update_write_addr_5__dout;
  wire update_write_addr_5__empty_n;
  wire update_write_addr_5__read;
  wire [64:0] update_write_addr_5__din;
  wire update_write_addr_5__full_n;
  wire update_write_addr_5__write;
  wire update_write_addr_5__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_addr_5__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_addr_5__rst__q2;
  wire [64:0] update_write_addr_6__dout;
  wire update_write_addr_6__empty_n;
  wire update_write_addr_6__read;
  wire [64:0] update_write_addr_6__din;
  wire update_write_addr_6__full_n;
  wire update_write_addr_6__write;
  wire update_write_addr_6__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_addr_6__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_addr_6__rst__q2;
  wire [64:0] update_write_addr_7__dout;
  wire update_write_addr_7__empty_n;
  wire update_write_addr_7__read;
  wire [64:0] update_write_addr_7__din;
  wire update_write_addr_7__full_n;
  wire update_write_addr_7__write;
  wire update_write_addr_7__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_addr_7__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_addr_7__rst__q2;
  wire [512:0] update_write_data_0__dout;
  wire update_write_data_0__empty_n;
  wire update_write_data_0__read;
  wire [512:0] update_write_data_0__din;
  wire update_write_data_0__full_n;
  wire update_write_data_0__write;
  wire update_write_data_0__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_data_0__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_data_0__rst__q2;
  wire [512:0] update_write_data_1__dout;
  wire update_write_data_1__empty_n;
  wire update_write_data_1__read;
  wire [512:0] update_write_data_1__din;
  wire update_write_data_1__full_n;
  wire update_write_data_1__write;
  wire update_write_data_1__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_data_1__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_data_1__rst__q2;
  wire [512:0] update_write_data_2__dout;
  wire update_write_data_2__empty_n;
  wire update_write_data_2__read;
  wire [512:0] update_write_data_2__din;
  wire update_write_data_2__full_n;
  wire update_write_data_2__write;
  wire update_write_data_2__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_data_2__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_data_2__rst__q2;
  wire [512:0] update_write_data_3__dout;
  wire update_write_data_3__empty_n;
  wire update_write_data_3__read;
  wire [512:0] update_write_data_3__din;
  wire update_write_data_3__full_n;
  wire update_write_data_3__write;
  wire update_write_data_3__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_data_3__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_data_3__rst__q2;
  wire [512:0] update_write_data_4__dout;
  wire update_write_data_4__empty_n;
  wire update_write_data_4__read;
  wire [512:0] update_write_data_4__din;
  wire update_write_data_4__full_n;
  wire update_write_data_4__write;
  wire update_write_data_4__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_data_4__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_data_4__rst__q2;
  wire [512:0] update_write_data_5__dout;
  wire update_write_data_5__empty_n;
  wire update_write_data_5__read;
  wire [512:0] update_write_data_5__din;
  wire update_write_data_5__full_n;
  wire update_write_data_5__write;
  wire update_write_data_5__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_data_5__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_data_5__rst__q2;
  wire [512:0] update_write_data_6__dout;
  wire update_write_data_6__empty_n;
  wire update_write_data_6__read;
  wire [512:0] update_write_data_6__din;
  wire update_write_data_6__full_n;
  wire update_write_data_6__write;
  wire update_write_data_6__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_data_6__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_data_6__rst__q2;
  wire [512:0] update_write_data_7__dout;
  wire update_write_data_7__empty_n;
  wire update_write_data_7__read;
  wire [512:0] update_write_data_7__din;
  wire update_write_data_7__full_n;
  wire update_write_data_7__write;
  wire update_write_data_7__rst__q0;
  (* dont_touch = "yes" *)
  reg update_write_data_7__rst__q1;
  (* dont_touch = "yes" *)
  reg update_write_data_7__rst__q2;
  wire [1024:0] vertex_mm2pe_r0_0__dout;
  wire vertex_mm2pe_r0_0__empty_n;
  wire vertex_mm2pe_r0_0__read;
  wire [1024:0] vertex_mm2pe_r0_0__din;
  wire vertex_mm2pe_r0_0__full_n;
  wire vertex_mm2pe_r0_0__write;
  wire vertex_mm2pe_r0_0__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r0_0__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r0_0__rst__q2;
  wire [1024:0] vertex_mm2pe_r0_1__dout;
  wire vertex_mm2pe_r0_1__empty_n;
  wire vertex_mm2pe_r0_1__read;
  wire [1024:0] vertex_mm2pe_r0_1__din;
  wire vertex_mm2pe_r0_1__full_n;
  wire vertex_mm2pe_r0_1__write;
  wire vertex_mm2pe_r0_1__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r0_1__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r0_1__rst__q2;
  wire [1024:0] vertex_mm2pe_r1_0__dout;
  wire vertex_mm2pe_r1_0__empty_n;
  wire vertex_mm2pe_r1_0__read;
  wire [1024:0] vertex_mm2pe_r1_0__din;
  wire vertex_mm2pe_r1_0__full_n;
  wire vertex_mm2pe_r1_0__write;
  wire vertex_mm2pe_r1_0__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r1_0__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r1_0__rst__q2;
  wire [1024:0] vertex_mm2pe_r1_1__dout;
  wire vertex_mm2pe_r1_1__empty_n;
  wire vertex_mm2pe_r1_1__read;
  wire [1024:0] vertex_mm2pe_r1_1__din;
  wire vertex_mm2pe_r1_1__full_n;
  wire vertex_mm2pe_r1_1__write;
  wire vertex_mm2pe_r1_1__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r1_1__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r1_1__rst__q2;
  wire [1024:0] vertex_mm2pe_r1_2__dout;
  wire vertex_mm2pe_r1_2__empty_n;
  wire vertex_mm2pe_r1_2__read;
  wire [1024:0] vertex_mm2pe_r1_2__din;
  wire vertex_mm2pe_r1_2__full_n;
  wire vertex_mm2pe_r1_2__write;
  wire vertex_mm2pe_r1_2__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r1_2__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r1_2__rst__q2;
  wire [1024:0] vertex_mm2pe_r1_3__dout;
  wire vertex_mm2pe_r1_3__empty_n;
  wire vertex_mm2pe_r1_3__read;
  wire [1024:0] vertex_mm2pe_r1_3__din;
  wire vertex_mm2pe_r1_3__full_n;
  wire vertex_mm2pe_r1_3__write;
  wire vertex_mm2pe_r1_3__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r1_3__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r1_3__rst__q2;
  wire [1024:0] vertex_mm2pe_r2_0__dout;
  wire vertex_mm2pe_r2_0__empty_n;
  wire vertex_mm2pe_r2_0__read;
  wire [1024:0] vertex_mm2pe_r2_0__din;
  wire vertex_mm2pe_r2_0__full_n;
  wire vertex_mm2pe_r2_0__write;
  wire vertex_mm2pe_r2_0__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r2_0__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r2_0__rst__q2;
  wire [1024:0] vertex_mm2pe_r2_1__dout;
  wire vertex_mm2pe_r2_1__empty_n;
  wire vertex_mm2pe_r2_1__read;
  wire [1024:0] vertex_mm2pe_r2_1__din;
  wire vertex_mm2pe_r2_1__full_n;
  wire vertex_mm2pe_r2_1__write;
  wire vertex_mm2pe_r2_1__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r2_1__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r2_1__rst__q2;
  wire [1024:0] vertex_mm2pe_r2_2__dout;
  wire vertex_mm2pe_r2_2__empty_n;
  wire vertex_mm2pe_r2_2__read;
  wire [1024:0] vertex_mm2pe_r2_2__din;
  wire vertex_mm2pe_r2_2__full_n;
  wire vertex_mm2pe_r2_2__write;
  wire vertex_mm2pe_r2_2__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r2_2__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r2_2__rst__q2;
  wire [1024:0] vertex_mm2pe_r2_3__dout;
  wire vertex_mm2pe_r2_3__empty_n;
  wire vertex_mm2pe_r2_3__read;
  wire [1024:0] vertex_mm2pe_r2_3__din;
  wire vertex_mm2pe_r2_3__full_n;
  wire vertex_mm2pe_r2_3__write;
  wire vertex_mm2pe_r2_3__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r2_3__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_mm2pe_r2_3__rst__q2;
  wire [1024:0] vertex_pe2mm_r0_0__dout;
  wire vertex_pe2mm_r0_0__empty_n;
  wire vertex_pe2mm_r0_0__read;
  wire [1024:0] vertex_pe2mm_r0_0__din;
  wire vertex_pe2mm_r0_0__full_n;
  wire vertex_pe2mm_r0_0__write;
  wire vertex_pe2mm_r0_0__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r0_0__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r0_0__rst__q2;
  wire [1024:0] vertex_pe2mm_r0_1__dout;
  wire vertex_pe2mm_r0_1__empty_n;
  wire vertex_pe2mm_r0_1__read;
  wire [1024:0] vertex_pe2mm_r0_1__din;
  wire vertex_pe2mm_r0_1__full_n;
  wire vertex_pe2mm_r0_1__write;
  wire vertex_pe2mm_r0_1__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r0_1__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r0_1__rst__q2;
  wire [1024:0] vertex_pe2mm_r1_0__dout;
  wire vertex_pe2mm_r1_0__empty_n;
  wire vertex_pe2mm_r1_0__read;
  wire [1024:0] vertex_pe2mm_r1_0__din;
  wire vertex_pe2mm_r1_0__full_n;
  wire vertex_pe2mm_r1_0__write;
  wire vertex_pe2mm_r1_0__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r1_0__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r1_0__rst__q2;
  wire [1024:0] vertex_pe2mm_r1_1__dout;
  wire vertex_pe2mm_r1_1__empty_n;
  wire vertex_pe2mm_r1_1__read;
  wire [1024:0] vertex_pe2mm_r1_1__din;
  wire vertex_pe2mm_r1_1__full_n;
  wire vertex_pe2mm_r1_1__write;
  wire vertex_pe2mm_r1_1__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r1_1__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r1_1__rst__q2;
  wire [1024:0] vertex_pe2mm_r1_2__dout;
  wire vertex_pe2mm_r1_2__empty_n;
  wire vertex_pe2mm_r1_2__read;
  wire [1024:0] vertex_pe2mm_r1_2__din;
  wire vertex_pe2mm_r1_2__full_n;
  wire vertex_pe2mm_r1_2__write;
  wire vertex_pe2mm_r1_2__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r1_2__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r1_2__rst__q2;
  wire [1024:0] vertex_pe2mm_r1_3__dout;
  wire vertex_pe2mm_r1_3__empty_n;
  wire vertex_pe2mm_r1_3__read;
  wire [1024:0] vertex_pe2mm_r1_3__din;
  wire vertex_pe2mm_r1_3__full_n;
  wire vertex_pe2mm_r1_3__write;
  wire vertex_pe2mm_r1_3__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r1_3__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r1_3__rst__q2;
  wire [1024:0] vertex_pe2mm_r2_0__dout;
  wire vertex_pe2mm_r2_0__empty_n;
  wire vertex_pe2mm_r2_0__read;
  wire [1024:0] vertex_pe2mm_r2_0__din;
  wire vertex_pe2mm_r2_0__full_n;
  wire vertex_pe2mm_r2_0__write;
  wire vertex_pe2mm_r2_0__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r2_0__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r2_0__rst__q2;
  wire [1024:0] vertex_pe2mm_r2_1__dout;
  wire vertex_pe2mm_r2_1__empty_n;
  wire vertex_pe2mm_r2_1__read;
  wire [1024:0] vertex_pe2mm_r2_1__din;
  wire vertex_pe2mm_r2_1__full_n;
  wire vertex_pe2mm_r2_1__write;
  wire vertex_pe2mm_r2_1__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r2_1__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r2_1__rst__q2;
  wire [1024:0] vertex_pe2mm_r2_2__dout;
  wire vertex_pe2mm_r2_2__empty_n;
  wire vertex_pe2mm_r2_2__read;
  wire [1024:0] vertex_pe2mm_r2_2__din;
  wire vertex_pe2mm_r2_2__full_n;
  wire vertex_pe2mm_r2_2__write;
  wire vertex_pe2mm_r2_2__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r2_2__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r2_2__rst__q2;
  wire [1024:0] vertex_pe2mm_r2_3__dout;
  wire vertex_pe2mm_r2_3__empty_n;
  wire vertex_pe2mm_r2_3__read;
  wire [1024:0] vertex_pe2mm_r2_3__din;
  wire vertex_pe2mm_r2_3__full_n;
  wire vertex_pe2mm_r2_3__write;
  wire vertex_pe2mm_r2_3__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r2_3__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_pe2mm_r2_3__rst__q2;
  wire [64:0] vertex_req_r0_0__dout;
  wire vertex_req_r0_0__empty_n;
  wire vertex_req_r0_0__read;
  wire [64:0] vertex_req_r0_0__din;
  wire vertex_req_r0_0__full_n;
  wire vertex_req_r0_0__write;
  wire vertex_req_r0_0__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r0_0__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r0_0__rst__q2;
  wire [64:0] vertex_req_r0_1__dout;
  wire vertex_req_r0_1__empty_n;
  wire vertex_req_r0_1__read;
  wire [64:0] vertex_req_r0_1__din;
  wire vertex_req_r0_1__full_n;
  wire vertex_req_r0_1__write;
  wire vertex_req_r0_1__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r0_1__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r0_1__rst__q2;
  wire [64:0] vertex_req_r1_0__dout;
  wire vertex_req_r1_0__empty_n;
  wire vertex_req_r1_0__read;
  wire [64:0] vertex_req_r1_0__din;
  wire vertex_req_r1_0__full_n;
  wire vertex_req_r1_0__write;
  wire vertex_req_r1_0__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r1_0__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r1_0__rst__q2;
  wire [64:0] vertex_req_r1_1__dout;
  wire vertex_req_r1_1__empty_n;
  wire vertex_req_r1_1__read;
  wire [64:0] vertex_req_r1_1__din;
  wire vertex_req_r1_1__full_n;
  wire vertex_req_r1_1__write;
  wire vertex_req_r1_1__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r1_1__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r1_1__rst__q2;
  wire [64:0] vertex_req_r1_2__dout;
  wire vertex_req_r1_2__empty_n;
  wire vertex_req_r1_2__read;
  wire [64:0] vertex_req_r1_2__din;
  wire vertex_req_r1_2__full_n;
  wire vertex_req_r1_2__write;
  wire vertex_req_r1_2__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r1_2__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r1_2__rst__q2;
  wire [64:0] vertex_req_r1_3__dout;
  wire vertex_req_r1_3__empty_n;
  wire vertex_req_r1_3__read;
  wire [64:0] vertex_req_r1_3__din;
  wire vertex_req_r1_3__full_n;
  wire vertex_req_r1_3__write;
  wire vertex_req_r1_3__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r1_3__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r1_3__rst__q2;
  wire [64:0] vertex_req_r2_0__dout;
  wire vertex_req_r2_0__empty_n;
  wire vertex_req_r2_0__read;
  wire [64:0] vertex_req_r2_0__din;
  wire vertex_req_r2_0__full_n;
  wire vertex_req_r2_0__write;
  wire vertex_req_r2_0__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r2_0__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r2_0__rst__q2;
  wire [64:0] vertex_req_r2_1__dout;
  wire vertex_req_r2_1__empty_n;
  wire vertex_req_r2_1__read;
  wire [64:0] vertex_req_r2_1__din;
  wire vertex_req_r2_1__full_n;
  wire vertex_req_r2_1__write;
  wire vertex_req_r2_1__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r2_1__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r2_1__rst__q2;
  wire [64:0] vertex_req_r2_2__dout;
  wire vertex_req_r2_2__empty_n;
  wire vertex_req_r2_2__read;
  wire [64:0] vertex_req_r2_2__din;
  wire vertex_req_r2_2__full_n;
  wire vertex_req_r2_2__write;
  wire vertex_req_r2_2__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r2_2__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r2_2__rst__q2;
  wire [64:0] vertex_req_r2_3__dout;
  wire vertex_req_r2_3__empty_n;
  wire vertex_req_r2_3__read;
  wire [64:0] vertex_req_r2_3__din;
  wire vertex_req_r2_3__full_n;
  wire vertex_req_r2_3__write;
  wire vertex_req_r2_3__rst__q0;
  (* dont_touch = "yes" *)
  reg vertex_req_r2_3__rst__q1;
  (* dont_touch = "yes" *)
  reg vertex_req_r2_3__rst__q2;
  wire [63:0] metadata__q0;
  (* dont_touch = "yes" *)
  reg [63:0] metadata__q1;
  (* dont_touch = "yes" *)
  reg [63:0] metadata__q2;
  wire [15:0] Control_0___num_partitions__q0;
  (* dont_touch = "yes" *)
  reg [15:0] Control_0___num_partitions__q1;
  (* dont_touch = "yes" *)
  reg [15:0] Control_0___num_partitions__q2;
  wire Control_0__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg Control_0__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg Control_0__ap_rst_n__q2;
  wire Control_0__is_done__q0;
  (* dont_touch = "yes" *)
  reg Control_0__is_done__q1;
  (* dont_touch = "yes" *)
  reg Control_0__is_done__q2;
  wire Control_0__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg Control_0__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg Control_0__ap_start_global__q2;
  wire Control_0__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg Control_0__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg Control_0__ap_done_global__q2;
  wire Control_0__ap_start;
  reg [1:0] Control_0__state;
  wire Control_0__ap_done;
  wire Control_0__ap_idle;
  wire Control_0__ap_ready;
  wire [63:0] edges_0__q0;
  (* dont_touch = "yes" *)
  reg [63:0] edges_0__q1;
  (* dont_touch = "yes" *)
  reg [63:0] edges_0__q2;
  wire [63:0] edges_0_read_addr__din;
  wire edges_0_read_addr__full_n;
  wire edges_0_read_addr__write;
  wire [511:0] edges_0_read_data__dout;
  wire edges_0_read_data__empty_n;
  wire edges_0_read_data__read;
  wire EdgeMem_0__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg EdgeMem_0__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg EdgeMem_0__ap_rst_n__q2;
  wire EdgeMem_0__ap_start;
  wire [63:0] edges_1__q0;
  (* dont_touch = "yes" *)
  reg [63:0] edges_1__q1;
  (* dont_touch = "yes" *)
  reg [63:0] edges_1__q2;
  wire [63:0] edges_1_read_addr__din;
  wire edges_1_read_addr__full_n;
  wire edges_1_read_addr__write;
  wire [511:0] edges_1_read_data__dout;
  wire edges_1_read_data__empty_n;
  wire edges_1_read_data__read;
  wire EdgeMem_1__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg EdgeMem_1__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg EdgeMem_1__ap_rst_n__q2;
  wire EdgeMem_1__ap_start;
  wire [63:0] edges_2__q0;
  (* dont_touch = "yes" *)
  reg [63:0] edges_2__q1;
  (* dont_touch = "yes" *)
  reg [63:0] edges_2__q2;
  wire [63:0] edges_2_read_addr__din;
  wire edges_2_read_addr__full_n;
  wire edges_2_read_addr__write;
  wire [511:0] edges_2_read_data__dout;
  wire edges_2_read_data__empty_n;
  wire edges_2_read_data__read;
  wire EdgeMem_2__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg EdgeMem_2__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg EdgeMem_2__ap_rst_n__q2;
  wire EdgeMem_2__ap_start;
  wire [63:0] edges_3__q0;
  (* dont_touch = "yes" *)
  reg [63:0] edges_3__q1;
  (* dont_touch = "yes" *)
  reg [63:0] edges_3__q2;
  wire [63:0] edges_3_read_addr__din;
  wire edges_3_read_addr__full_n;
  wire edges_3_read_addr__write;
  wire [511:0] edges_3_read_data__dout;
  wire edges_3_read_data__empty_n;
  wire edges_3_read_data__read;
  wire EdgeMem_3__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg EdgeMem_3__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg EdgeMem_3__ap_rst_n__q2;
  wire EdgeMem_3__ap_start;
  wire [63:0] edges_4__q0;
  (* dont_touch = "yes" *)
  reg [63:0] edges_4__q1;
  (* dont_touch = "yes" *)
  reg [63:0] edges_4__q2;
  wire [63:0] edges_4_read_addr__din;
  wire edges_4_read_addr__full_n;
  wire edges_4_read_addr__write;
  wire [511:0] edges_4_read_data__dout;
  wire edges_4_read_data__empty_n;
  wire edges_4_read_data__read;
  wire EdgeMem_4__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg EdgeMem_4__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg EdgeMem_4__ap_rst_n__q2;
  wire EdgeMem_4__ap_start;
  wire [63:0] edges_5__q0;
  (* dont_touch = "yes" *)
  reg [63:0] edges_5__q1;
  (* dont_touch = "yes" *)
  reg [63:0] edges_5__q2;
  wire [63:0] edges_5_read_addr__din;
  wire edges_5_read_addr__full_n;
  wire edges_5_read_addr__write;
  wire [511:0] edges_5_read_data__dout;
  wire edges_5_read_data__empty_n;
  wire edges_5_read_data__read;
  wire EdgeMem_5__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg EdgeMem_5__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg EdgeMem_5__ap_rst_n__q2;
  wire EdgeMem_5__ap_start;
  wire [63:0] edges_6__q0;
  (* dont_touch = "yes" *)
  reg [63:0] edges_6__q1;
  (* dont_touch = "yes" *)
  reg [63:0] edges_6__q2;
  wire [63:0] edges_6_read_addr__din;
  wire edges_6_read_addr__full_n;
  wire edges_6_read_addr__write;
  wire [511:0] edges_6_read_data__dout;
  wire edges_6_read_data__empty_n;
  wire edges_6_read_data__read;
  wire EdgeMem_6__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg EdgeMem_6__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg EdgeMem_6__ap_rst_n__q2;
  wire EdgeMem_6__ap_start;
  wire [63:0] edges_7__q0;
  (* dont_touch = "yes" *)
  reg [63:0] edges_7__q1;
  (* dont_touch = "yes" *)
  reg [63:0] edges_7__q2;
  wire [63:0] edges_7_read_addr__din;
  wire edges_7_read_addr__full_n;
  wire edges_7_read_addr__write;
  wire [511:0] edges_7_read_data__dout;
  wire edges_7_read_data__empty_n;
  wire edges_7_read_data__read;
  wire EdgeMem_7__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg EdgeMem_7__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg EdgeMem_7__ap_rst_n__q2;
  wire EdgeMem_7__ap_start;
  wire ProcElem_0__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_0__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_0__ap_rst_n__q2;
  wire ProcElem_0__is_done__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_0__is_done__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_0__is_done__q2;
  wire ProcElem_0__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_0__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_0__ap_start_global__q2;
  wire ProcElem_0__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_0__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_0__ap_done_global__q2;
  wire ProcElem_0__ap_start;
  reg [1:0] ProcElem_0__state;
  wire ProcElem_0__ap_done;
  wire ProcElem_0__ap_idle;
  wire ProcElem_0__ap_ready;
  wire ProcElem_1__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_1__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_1__ap_rst_n__q2;
  wire ProcElem_1__is_done__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_1__is_done__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_1__is_done__q2;
  wire ProcElem_1__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_1__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_1__ap_start_global__q2;
  wire ProcElem_1__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_1__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_1__ap_done_global__q2;
  wire ProcElem_1__ap_start;
  reg [1:0] ProcElem_1__state;
  wire ProcElem_1__ap_done;
  wire ProcElem_1__ap_idle;
  wire ProcElem_1__ap_ready;
  wire ProcElem_2__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_2__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_2__ap_rst_n__q2;
  wire ProcElem_2__is_done__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_2__is_done__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_2__is_done__q2;
  wire ProcElem_2__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_2__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_2__ap_start_global__q2;
  wire ProcElem_2__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_2__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_2__ap_done_global__q2;
  wire ProcElem_2__ap_start;
  reg [1:0] ProcElem_2__state;
  wire ProcElem_2__ap_done;
  wire ProcElem_2__ap_idle;
  wire ProcElem_2__ap_ready;
  wire ProcElem_3__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_3__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_3__ap_rst_n__q2;
  wire ProcElem_3__is_done__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_3__is_done__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_3__is_done__q2;
  wire ProcElem_3__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_3__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_3__ap_start_global__q2;
  wire ProcElem_3__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_3__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_3__ap_done_global__q2;
  wire ProcElem_3__ap_start;
  reg [1:0] ProcElem_3__state;
  wire ProcElem_3__ap_done;
  wire ProcElem_3__ap_idle;
  wire ProcElem_3__ap_ready;
  wire ProcElem_4__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_4__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_4__ap_rst_n__q2;
  wire ProcElem_4__is_done__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_4__is_done__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_4__is_done__q2;
  wire ProcElem_4__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_4__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_4__ap_start_global__q2;
  wire ProcElem_4__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_4__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_4__ap_done_global__q2;
  wire ProcElem_4__ap_start;
  reg [1:0] ProcElem_4__state;
  wire ProcElem_4__ap_done;
  wire ProcElem_4__ap_idle;
  wire ProcElem_4__ap_ready;
  wire ProcElem_5__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_5__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_5__ap_rst_n__q2;
  wire ProcElem_5__is_done__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_5__is_done__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_5__is_done__q2;
  wire ProcElem_5__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_5__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_5__ap_start_global__q2;
  wire ProcElem_5__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_5__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_5__ap_done_global__q2;
  wire ProcElem_5__ap_start;
  reg [1:0] ProcElem_5__state;
  wire ProcElem_5__ap_done;
  wire ProcElem_5__ap_idle;
  wire ProcElem_5__ap_ready;
  wire ProcElem_6__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_6__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_6__ap_rst_n__q2;
  wire ProcElem_6__is_done__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_6__is_done__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_6__is_done__q2;
  wire ProcElem_6__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_6__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_6__ap_start_global__q2;
  wire ProcElem_6__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_6__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_6__ap_done_global__q2;
  wire ProcElem_6__ap_start;
  reg [1:0] ProcElem_6__state;
  wire ProcElem_6__ap_done;
  wire ProcElem_6__ap_idle;
  wire ProcElem_6__ap_ready;
  wire ProcElem_7__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_7__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_7__ap_rst_n__q2;
  wire ProcElem_7__is_done__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_7__is_done__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_7__is_done__q2;
  wire ProcElem_7__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_7__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_7__ap_start_global__q2;
  wire ProcElem_7__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg ProcElem_7__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg ProcElem_7__ap_done_global__q2;
  wire ProcElem_7__ap_start;
  reg [1:0] ProcElem_7__state;
  wire ProcElem_7__ap_done;
  wire ProcElem_7__ap_idle;
  wire ProcElem_7__ap_ready;
  wire [15:0] UpdateHandler_0___num_partitions__q0;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_0___num_partitions__q1;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_0___num_partitions__q2;
  wire UpdateHandler_0__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_0__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_0__ap_rst_n__q2;
  wire UpdateHandler_0__is_done__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_0__is_done__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_0__is_done__q2;
  wire UpdateHandler_0__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_0__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_0__ap_start_global__q2;
  wire UpdateHandler_0__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_0__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_0__ap_done_global__q2;
  wire UpdateHandler_0__ap_start;
  reg [1:0] UpdateHandler_0__state;
  wire UpdateHandler_0__ap_done;
  wire UpdateHandler_0__ap_idle;
  wire UpdateHandler_0__ap_ready;
  wire [15:0] UpdateHandler_1___num_partitions__q0;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_1___num_partitions__q1;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_1___num_partitions__q2;
  wire UpdateHandler_1__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_1__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_1__ap_rst_n__q2;
  wire UpdateHandler_1__is_done__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_1__is_done__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_1__is_done__q2;
  wire UpdateHandler_1__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_1__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_1__ap_start_global__q2;
  wire UpdateHandler_1__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_1__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_1__ap_done_global__q2;
  wire UpdateHandler_1__ap_start;
  reg [1:0] UpdateHandler_1__state;
  wire UpdateHandler_1__ap_done;
  wire UpdateHandler_1__ap_idle;
  wire UpdateHandler_1__ap_ready;
  wire [15:0] UpdateHandler_2___num_partitions__q0;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_2___num_partitions__q1;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_2___num_partitions__q2;
  wire UpdateHandler_2__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_2__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_2__ap_rst_n__q2;
  wire UpdateHandler_2__is_done__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_2__is_done__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_2__is_done__q2;
  wire UpdateHandler_2__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_2__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_2__ap_start_global__q2;
  wire UpdateHandler_2__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_2__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_2__ap_done_global__q2;
  wire UpdateHandler_2__ap_start;
  reg [1:0] UpdateHandler_2__state;
  wire UpdateHandler_2__ap_done;
  wire UpdateHandler_2__ap_idle;
  wire UpdateHandler_2__ap_ready;
  wire [15:0] UpdateHandler_3___num_partitions__q0;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_3___num_partitions__q1;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_3___num_partitions__q2;
  wire UpdateHandler_3__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_3__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_3__ap_rst_n__q2;
  wire UpdateHandler_3__is_done__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_3__is_done__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_3__is_done__q2;
  wire UpdateHandler_3__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_3__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_3__ap_start_global__q2;
  wire UpdateHandler_3__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_3__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_3__ap_done_global__q2;
  wire UpdateHandler_3__ap_start;
  reg [1:0] UpdateHandler_3__state;
  wire UpdateHandler_3__ap_done;
  wire UpdateHandler_3__ap_idle;
  wire UpdateHandler_3__ap_ready;
  wire [15:0] UpdateHandler_4___num_partitions__q0;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_4___num_partitions__q1;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_4___num_partitions__q2;
  wire UpdateHandler_4__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_4__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_4__ap_rst_n__q2;
  wire UpdateHandler_4__is_done__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_4__is_done__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_4__is_done__q2;
  wire UpdateHandler_4__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_4__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_4__ap_start_global__q2;
  wire UpdateHandler_4__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_4__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_4__ap_done_global__q2;
  wire UpdateHandler_4__ap_start;
  reg [1:0] UpdateHandler_4__state;
  wire UpdateHandler_4__ap_done;
  wire UpdateHandler_4__ap_idle;
  wire UpdateHandler_4__ap_ready;
  wire [15:0] UpdateHandler_5___num_partitions__q0;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_5___num_partitions__q1;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_5___num_partitions__q2;
  wire UpdateHandler_5__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_5__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_5__ap_rst_n__q2;
  wire UpdateHandler_5__is_done__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_5__is_done__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_5__is_done__q2;
  wire UpdateHandler_5__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_5__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_5__ap_start_global__q2;
  wire UpdateHandler_5__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_5__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_5__ap_done_global__q2;
  wire UpdateHandler_5__ap_start;
  reg [1:0] UpdateHandler_5__state;
  wire UpdateHandler_5__ap_done;
  wire UpdateHandler_5__ap_idle;
  wire UpdateHandler_5__ap_ready;
  wire [15:0] UpdateHandler_6___num_partitions__q0;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_6___num_partitions__q1;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_6___num_partitions__q2;
  wire UpdateHandler_6__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_6__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_6__ap_rst_n__q2;
  wire UpdateHandler_6__is_done__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_6__is_done__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_6__is_done__q2;
  wire UpdateHandler_6__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_6__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_6__ap_start_global__q2;
  wire UpdateHandler_6__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_6__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_6__ap_done_global__q2;
  wire UpdateHandler_6__ap_start;
  reg [1:0] UpdateHandler_6__state;
  wire UpdateHandler_6__ap_done;
  wire UpdateHandler_6__ap_idle;
  wire UpdateHandler_6__ap_ready;
  wire [15:0] UpdateHandler_7___num_partitions__q0;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_7___num_partitions__q1;
  (* dont_touch = "yes" *)
  reg [15:0] UpdateHandler_7___num_partitions__q2;
  wire UpdateHandler_7__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_7__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_7__ap_rst_n__q2;
  wire UpdateHandler_7__is_done__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_7__is_done__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_7__is_done__q2;
  wire UpdateHandler_7__ap_start_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_7__ap_start_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_7__ap_start_global__q2;
  wire UpdateHandler_7__ap_done_global__q0;
  (* dont_touch = "yes" *)
  reg UpdateHandler_7__ap_done_global__q1;
  (* dont_touch = "yes" *)
  reg UpdateHandler_7__ap_done_global__q2;
  wire UpdateHandler_7__ap_start;
  reg [1:0] UpdateHandler_7__state;
  wire UpdateHandler_7__ap_done;
  wire UpdateHandler_7__ap_idle;
  wire UpdateHandler_7__ap_ready;
  wire [63:0] updates_0__q0;
  (* dont_touch = "yes" *)
  reg [63:0] updates_0__q1;
  (* dont_touch = "yes" *)
  reg [63:0] updates_0__q2;
  wire [63:0] updates_0_read_addr__din;
  wire updates_0_read_addr__full_n;
  wire updates_0_read_addr__write;
  wire [511:0] updates_0_read_data__dout;
  wire updates_0_read_data__empty_n;
  wire updates_0_read_data__read;
  wire [63:0] updates_0_write_addr__din;
  wire updates_0_write_addr__full_n;
  wire updates_0_write_addr__write;
  wire [511:0] updates_0_write_data__din;
  wire updates_0_write_data__full_n;
  wire updates_0_write_data__write;
  wire UpdateMem_0__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateMem_0__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateMem_0__ap_rst_n__q2;
  wire UpdateMem_0__ap_start;
  wire [63:0] updates_1__q0;
  (* dont_touch = "yes" *)
  reg [63:0] updates_1__q1;
  (* dont_touch = "yes" *)
  reg [63:0] updates_1__q2;
  wire [63:0] updates_1_read_addr__din;
  wire updates_1_read_addr__full_n;
  wire updates_1_read_addr__write;
  wire [511:0] updates_1_read_data__dout;
  wire updates_1_read_data__empty_n;
  wire updates_1_read_data__read;
  wire [63:0] updates_1_write_addr__din;
  wire updates_1_write_addr__full_n;
  wire updates_1_write_addr__write;
  wire [511:0] updates_1_write_data__din;
  wire updates_1_write_data__full_n;
  wire updates_1_write_data__write;
  wire UpdateMem_1__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateMem_1__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateMem_1__ap_rst_n__q2;
  wire UpdateMem_1__ap_start;
  wire [63:0] updates_2__q0;
  (* dont_touch = "yes" *)
  reg [63:0] updates_2__q1;
  (* dont_touch = "yes" *)
  reg [63:0] updates_2__q2;
  wire [63:0] updates_2_read_addr__din;
  wire updates_2_read_addr__full_n;
  wire updates_2_read_addr__write;
  wire [511:0] updates_2_read_data__dout;
  wire updates_2_read_data__empty_n;
  wire updates_2_read_data__read;
  wire [63:0] updates_2_write_addr__din;
  wire updates_2_write_addr__full_n;
  wire updates_2_write_addr__write;
  wire [511:0] updates_2_write_data__din;
  wire updates_2_write_data__full_n;
  wire updates_2_write_data__write;
  wire UpdateMem_2__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateMem_2__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateMem_2__ap_rst_n__q2;
  wire UpdateMem_2__ap_start;
  wire [63:0] updates_3__q0;
  (* dont_touch = "yes" *)
  reg [63:0] updates_3__q1;
  (* dont_touch = "yes" *)
  reg [63:0] updates_3__q2;
  wire [63:0] updates_3_read_addr__din;
  wire updates_3_read_addr__full_n;
  wire updates_3_read_addr__write;
  wire [511:0] updates_3_read_data__dout;
  wire updates_3_read_data__empty_n;
  wire updates_3_read_data__read;
  wire [63:0] updates_3_write_addr__din;
  wire updates_3_write_addr__full_n;
  wire updates_3_write_addr__write;
  wire [511:0] updates_3_write_data__din;
  wire updates_3_write_data__full_n;
  wire updates_3_write_data__write;
  wire UpdateMem_3__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateMem_3__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateMem_3__ap_rst_n__q2;
  wire UpdateMem_3__ap_start;
  wire [63:0] updates_4__q0;
  (* dont_touch = "yes" *)
  reg [63:0] updates_4__q1;
  (* dont_touch = "yes" *)
  reg [63:0] updates_4__q2;
  wire [63:0] updates_4_read_addr__din;
  wire updates_4_read_addr__full_n;
  wire updates_4_read_addr__write;
  wire [511:0] updates_4_read_data__dout;
  wire updates_4_read_data__empty_n;
  wire updates_4_read_data__read;
  wire [63:0] updates_4_write_addr__din;
  wire updates_4_write_addr__full_n;
  wire updates_4_write_addr__write;
  wire [511:0] updates_4_write_data__din;
  wire updates_4_write_data__full_n;
  wire updates_4_write_data__write;
  wire UpdateMem_4__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateMem_4__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateMem_4__ap_rst_n__q2;
  wire UpdateMem_4__ap_start;
  wire [63:0] updates_5__q0;
  (* dont_touch = "yes" *)
  reg [63:0] updates_5__q1;
  (* dont_touch = "yes" *)
  reg [63:0] updates_5__q2;
  wire [63:0] updates_5_read_addr__din;
  wire updates_5_read_addr__full_n;
  wire updates_5_read_addr__write;
  wire [511:0] updates_5_read_data__dout;
  wire updates_5_read_data__empty_n;
  wire updates_5_read_data__read;
  wire [63:0] updates_5_write_addr__din;
  wire updates_5_write_addr__full_n;
  wire updates_5_write_addr__write;
  wire [511:0] updates_5_write_data__din;
  wire updates_5_write_data__full_n;
  wire updates_5_write_data__write;
  wire UpdateMem_5__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateMem_5__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateMem_5__ap_rst_n__q2;
  wire UpdateMem_5__ap_start;
  wire [63:0] updates_6__q0;
  (* dont_touch = "yes" *)
  reg [63:0] updates_6__q1;
  (* dont_touch = "yes" *)
  reg [63:0] updates_6__q2;
  wire [63:0] updates_6_read_addr__din;
  wire updates_6_read_addr__full_n;
  wire updates_6_read_addr__write;
  wire [511:0] updates_6_read_data__dout;
  wire updates_6_read_data__empty_n;
  wire updates_6_read_data__read;
  wire [63:0] updates_6_write_addr__din;
  wire updates_6_write_addr__full_n;
  wire updates_6_write_addr__write;
  wire [511:0] updates_6_write_data__din;
  wire updates_6_write_data__full_n;
  wire updates_6_write_data__write;
  wire UpdateMem_6__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateMem_6__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateMem_6__ap_rst_n__q2;
  wire UpdateMem_6__ap_start;
  wire [63:0] updates_7__q0;
  (* dont_touch = "yes" *)
  reg [63:0] updates_7__q1;
  (* dont_touch = "yes" *)
  reg [63:0] updates_7__q2;
  wire [63:0] updates_7_read_addr__din;
  wire updates_7_read_addr__full_n;
  wire updates_7_read_addr__write;
  wire [511:0] updates_7_read_data__dout;
  wire updates_7_read_data__empty_n;
  wire updates_7_read_data__read;
  wire [63:0] updates_7_write_addr__din;
  wire updates_7_write_addr__full_n;
  wire updates_7_write_addr__write;
  wire [511:0] updates_7_write_data__din;
  wire updates_7_write_data__full_n;
  wire updates_7_write_data__write;
  wire UpdateMem_7__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg UpdateMem_7__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg UpdateMem_7__ap_rst_n__q2;
  wire UpdateMem_7__ap_start;
  wire [63:0] degrees__q0;
  (* dont_touch = "yes" *)
  reg [63:0] degrees__q1;
  (* dont_touch = "yes" *)
  reg [63:0] degrees__q2;
  wire [63:0] degrees_read_addr__din;
  wire degrees_read_addr__full_n;
  wire degrees_read_addr__write;
  wire [511:0] degrees_read_data__dout;
  wire degrees_read_data__empty_n;
  wire degrees_read_data__read;
  wire [63:0] rankings__q0;
  (* dont_touch = "yes" *)
  reg [63:0] rankings__q1;
  (* dont_touch = "yes" *)
  reg [63:0] rankings__q2;
  wire [63:0] rankings_read_addr__din;
  wire rankings_read_addr__full_n;
  wire rankings_read_addr__write;
  wire [511:0] rankings_read_data__dout;
  wire rankings_read_data__empty_n;
  wire rankings_read_data__read;
  wire [63:0] rankings_write_addr__din;
  wire rankings_write_addr__full_n;
  wire rankings_write_addr__write;
  wire [511:0] rankings_write_data__din;
  wire rankings_write_data__full_n;
  wire rankings_write_data__write;
  wire [63:0] tmps__q0;
  (* dont_touch = "yes" *)
  reg [63:0] tmps__q1;
  (* dont_touch = "yes" *)
  reg [63:0] tmps__q2;
  wire [63:0] tmps_read_addr__din;
  wire tmps_read_addr__full_n;
  wire tmps_read_addr__write;
  wire [511:0] tmps_read_data__dout;
  wire tmps_read_data__empty_n;
  wire tmps_read_data__read;
  wire [63:0] tmps_write_addr__din;
  wire tmps_write_addr__full_n;
  wire tmps_write_addr__write;
  wire [511:0] tmps_write_data__din;
  wire tmps_write_data__full_n;
  wire tmps_write_data__write;
  wire VertexMem_0__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg VertexMem_0__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg VertexMem_0__ap_rst_n__q2;
  wire VertexMem_0__ap_start;
  wire VertexRouterR1_0__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg VertexRouterR1_0__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg VertexRouterR1_0__ap_rst_n__q2;
  wire VertexRouterR1_0__ap_start;
  wire VertexRouterR2_0__ap_rst_n__q0;
  (* dont_touch = "yes" *)
  reg VertexRouterR2_0__ap_rst_n__q1;
  (* dont_touch = "yes" *)
  reg VertexRouterR2_0__ap_rst_n__q2;
  wire VertexRouterR2_0__ap_start;
  wire edges_0__rst__q0;
  (* dont_touch = "yes" *)
  reg edges_0__rst__q1;
  (* dont_touch = "yes" *)
  reg edges_0__rst__q2;
  wire edges_1__rst__q0;
  (* dont_touch = "yes" *)
  reg edges_1__rst__q1;
  (* dont_touch = "yes" *)
  reg edges_1__rst__q2;
  wire edges_2__rst__q0;
  (* dont_touch = "yes" *)
  reg edges_2__rst__q1;
  (* dont_touch = "yes" *)
  reg edges_2__rst__q2;
  wire edges_3__rst__q0;
  (* dont_touch = "yes" *)
  reg edges_3__rst__q1;
  (* dont_touch = "yes" *)
  reg edges_3__rst__q2;
  wire edges_4__rst__q0;
  (* dont_touch = "yes" *)
  reg edges_4__rst__q1;
  (* dont_touch = "yes" *)
  reg edges_4__rst__q2;
  wire edges_5__rst__q0;
  (* dont_touch = "yes" *)
  reg edges_5__rst__q1;
  (* dont_touch = "yes" *)
  reg edges_5__rst__q2;
  wire edges_6__rst__q0;
  (* dont_touch = "yes" *)
  reg edges_6__rst__q1;
  (* dont_touch = "yes" *)
  reg edges_6__rst__q2;
  wire edges_7__rst__q0;
  (* dont_touch = "yes" *)
  reg edges_7__rst__q1;
  (* dont_touch = "yes" *)
  reg edges_7__rst__q2;
  wire updates_0__rst__q0;
  (* dont_touch = "yes" *)
  reg updates_0__rst__q1;
  (* dont_touch = "yes" *)
  reg updates_0__rst__q2;
  wire updates_1__rst__q0;
  (* dont_touch = "yes" *)
  reg updates_1__rst__q1;
  (* dont_touch = "yes" *)
  reg updates_1__rst__q2;
  wire updates_2__rst__q0;
  (* dont_touch = "yes" *)
  reg updates_2__rst__q1;
  (* dont_touch = "yes" *)
  reg updates_2__rst__q2;
  wire updates_3__rst__q0;
  (* dont_touch = "yes" *)
  reg updates_3__rst__q1;
  (* dont_touch = "yes" *)
  reg updates_3__rst__q2;
  wire updates_4__rst__q0;
  (* dont_touch = "yes" *)
  reg updates_4__rst__q1;
  (* dont_touch = "yes" *)
  reg updates_4__rst__q2;
  wire updates_5__rst__q0;
  (* dont_touch = "yes" *)
  reg updates_5__rst__q1;
  (* dont_touch = "yes" *)
  reg updates_5__rst__q2;
  wire updates_6__rst__q0;
  (* dont_touch = "yes" *)
  reg updates_6__rst__q1;
  (* dont_touch = "yes" *)
  reg updates_6__rst__q2;
  wire updates_7__rst__q0;
  (* dont_touch = "yes" *)
  reg updates_7__rst__q1;
  (* dont_touch = "yes" *)
  reg updates_7__rst__q2;
  wire degrees__rst__q0;
  (* dont_touch = "yes" *)
  reg degrees__rst__q1;
  (* dont_touch = "yes" *)
  reg degrees__rst__q2;
  wire rankings__rst__q0;
  (* dont_touch = "yes" *)
  reg rankings__rst__q1;
  (* dont_touch = "yes" *)
  reg rankings__rst__q2;
  wire tmps__rst__q0;
  (* dont_touch = "yes" *)
  reg tmps__rst__q1;
  (* dont_touch = "yes" *)
  reg tmps__rst__q2;
  reg [1:0] tlp_state;
  reg [0:0] countdown;
  wire ap_start__q0;
  (* dont_touch = "yes" *)
  reg ap_start__q1;
  (* dont_touch = "yes" *)
  reg ap_start__q2;
  wire ap_done__q0;
  (* dont_touch = "yes" *)
  reg ap_done__q1;
  (* dont_touch = "yes" *)
  reg ap_done__q2;

  PageRank_PageRank_control_s_axi
  #(
    .C_S_AXI_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_S_AXI_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH)
  )
  PageRank_control_s_axi_U
  (
    .AWVALID(s_axi_control_AWVALID),
    .AWREADY(s_axi_control_AWREADY),
    .AWADDR(s_axi_control_AWADDR),
    .WVALID(s_axi_control_WVALID),
    .WREADY(s_axi_control_WREADY),
    .WDATA(s_axi_control_WDATA),
    .WSTRB(s_axi_control_WSTRB),
    .ARVALID(s_axi_control_ARVALID),
    .ARREADY(s_axi_control_ARREADY),
    .ARADDR(s_axi_control_ARADDR),
    .RVALID(s_axi_control_RVALID),
    .RREADY(s_axi_control_RREADY),
    .RDATA(s_axi_control_RDATA),
    .RRESP(s_axi_control_RRESP),
    .BVALID(s_axi_control_BVALID),
    .BREADY(s_axi_control_BREADY),
    .BRESP(s_axi_control_BRESP),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .ap_start(ap_start),
    .interrupt(interrupt),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .num_partitions(num_partitions),
    .metadata(metadata),
    .degrees(degrees),
    .rankings(rankings),
    .tmps(tmps),
    .edges_0(edges_0),
    .edges_1(edges_1),
    .edges_2(edges_2),
    .edges_3(edges_3),
    .edges_4(edges_4),
    .edges_5(edges_5),
    .edges_6(edges_6),
    .edges_7(edges_7),
    .updates_0(updates_0),
    .updates_1(updates_1),
    .updates_2(updates_2),
    .updates_3(updates_3),
    .updates_4(updates_4),
    .updates_5(updates_5),
    .updates_6(updates_6),
    .updates_7(updates_7)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_req_0
  (
    .clk(ap_clk),
    .reset(edge_req_0__rst__q2),
    .if_dout(edge_req_0__dout),
    .if_empty_n(edge_req_0__empty_n),
    .if_read(edge_req_0__read),
    .if_read_ce(1'b1),
    .if_din(edge_req_0__din),
    .if_full_n(edge_req_0__full_n),
    .if_write(edge_req_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_req_1
  (
    .clk(ap_clk),
    .reset(edge_req_1__rst__q2),
    .if_dout(edge_req_1__dout),
    .if_empty_n(edge_req_1__empty_n),
    .if_read(edge_req_1__read),
    .if_read_ce(1'b1),
    .if_din(edge_req_1__din),
    .if_full_n(edge_req_1__full_n),
    .if_write(edge_req_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_req_2
  (
    .clk(ap_clk),
    .reset(edge_req_2__rst__q2),
    .if_dout(edge_req_2__dout),
    .if_empty_n(edge_req_2__empty_n),
    .if_read(edge_req_2__read),
    .if_read_ce(1'b1),
    .if_din(edge_req_2__din),
    .if_full_n(edge_req_2__full_n),
    .if_write(edge_req_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_req_3
  (
    .clk(ap_clk),
    .reset(edge_req_3__rst__q2),
    .if_dout(edge_req_3__dout),
    .if_empty_n(edge_req_3__empty_n),
    .if_read(edge_req_3__read),
    .if_read_ce(1'b1),
    .if_din(edge_req_3__din),
    .if_full_n(edge_req_3__full_n),
    .if_write(edge_req_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_req_4
  (
    .clk(ap_clk),
    .reset(edge_req_4__rst__q2),
    .if_dout(edge_req_4__dout),
    .if_empty_n(edge_req_4__empty_n),
    .if_read(edge_req_4__read),
    .if_read_ce(1'b1),
    .if_din(edge_req_4__din),
    .if_full_n(edge_req_4__full_n),
    .if_write(edge_req_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_req_5
  (
    .clk(ap_clk),
    .reset(edge_req_5__rst__q2),
    .if_dout(edge_req_5__dout),
    .if_empty_n(edge_req_5__empty_n),
    .if_read(edge_req_5__read),
    .if_read_ce(1'b1),
    .if_din(edge_req_5__din),
    .if_full_n(edge_req_5__full_n),
    .if_write(edge_req_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_req_6
  (
    .clk(ap_clk),
    .reset(edge_req_6__rst__q2),
    .if_dout(edge_req_6__dout),
    .if_empty_n(edge_req_6__empty_n),
    .if_read(edge_req_6__read),
    .if_read_ce(1'b1),
    .if_din(edge_req_6__din),
    .if_full_n(edge_req_6__full_n),
    .if_write(edge_req_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_req_7
  (
    .clk(ap_clk),
    .reset(edge_req_7__rst__q2),
    .if_dout(edge_req_7__dout),
    .if_empty_n(edge_req_7__empty_n),
    .if_read(edge_req_7__read),
    .if_read_ce(1'b1),
    .if_din(edge_req_7__din),
    .if_full_n(edge_req_7__full_n),
    .if_write(edge_req_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_resp_0
  (
    .clk(ap_clk),
    .reset(edge_resp_0__rst__q2),
    .if_dout(edge_resp_0__dout),
    .if_empty_n(edge_resp_0__empty_n),
    .if_read(edge_resp_0__read),
    .if_read_ce(1'b1),
    .if_din(edge_resp_0__din),
    .if_full_n(edge_resp_0__full_n),
    .if_write(edge_resp_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_resp_1
  (
    .clk(ap_clk),
    .reset(edge_resp_1__rst__q2),
    .if_dout(edge_resp_1__dout),
    .if_empty_n(edge_resp_1__empty_n),
    .if_read(edge_resp_1__read),
    .if_read_ce(1'b1),
    .if_din(edge_resp_1__din),
    .if_full_n(edge_resp_1__full_n),
    .if_write(edge_resp_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_resp_2
  (
    .clk(ap_clk),
    .reset(edge_resp_2__rst__q2),
    .if_dout(edge_resp_2__dout),
    .if_empty_n(edge_resp_2__empty_n),
    .if_read(edge_resp_2__read),
    .if_read_ce(1'b1),
    .if_din(edge_resp_2__din),
    .if_full_n(edge_resp_2__full_n),
    .if_write(edge_resp_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_resp_3
  (
    .clk(ap_clk),
    .reset(edge_resp_3__rst__q2),
    .if_dout(edge_resp_3__dout),
    .if_empty_n(edge_resp_3__empty_n),
    .if_read(edge_resp_3__read),
    .if_read_ce(1'b1),
    .if_din(edge_resp_3__din),
    .if_full_n(edge_resp_3__full_n),
    .if_write(edge_resp_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_resp_4
  (
    .clk(ap_clk),
    .reset(edge_resp_4__rst__q2),
    .if_dout(edge_resp_4__dout),
    .if_empty_n(edge_resp_4__empty_n),
    .if_read(edge_resp_4__read),
    .if_read_ce(1'b1),
    .if_din(edge_resp_4__din),
    .if_full_n(edge_resp_4__full_n),
    .if_write(edge_resp_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_resp_5
  (
    .clk(ap_clk),
    .reset(edge_resp_5__rst__q2),
    .if_dout(edge_resp_5__dout),
    .if_empty_n(edge_resp_5__empty_n),
    .if_read(edge_resp_5__read),
    .if_read_ce(1'b1),
    .if_din(edge_resp_5__din),
    .if_full_n(edge_resp_5__full_n),
    .if_write(edge_resp_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_resp_6
  (
    .clk(ap_clk),
    .reset(edge_resp_6__rst__q2),
    .if_dout(edge_resp_6__dout),
    .if_empty_n(edge_resp_6__empty_n),
    .if_read(edge_resp_6__read),
    .if_read_ce(1'b1),
    .if_din(edge_resp_6__din),
    .if_full_n(edge_resp_6__full_n),
    .if_write(edge_resp_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  edge_resp_7
  (
    .clk(ap_clk),
    .reset(edge_resp_7__rst__q2),
    .if_dout(edge_resp_7__dout),
    .if_empty_n(edge_resp_7__empty_n),
    .if_read(edge_resp_7__read),
    .if_read_ce(1'b1),
    .if_din(edge_resp_7__din),
    .if_full_n(edge_resp_7__full_n),
    .if_write(edge_resp_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(49),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  num_updates_0
  (
    .clk(ap_clk),
    .reset(num_updates_0__rst__q2),
    .if_dout(num_updates_0__dout),
    .if_empty_n(num_updates_0__empty_n),
    .if_read(num_updates_0__read),
    .if_read_ce(1'b1),
    .if_din(num_updates_0__din),
    .if_full_n(num_updates_0__full_n),
    .if_write(num_updates_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(49),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  num_updates_1
  (
    .clk(ap_clk),
    .reset(num_updates_1__rst__q2),
    .if_dout(num_updates_1__dout),
    .if_empty_n(num_updates_1__empty_n),
    .if_read(num_updates_1__read),
    .if_read_ce(1'b1),
    .if_din(num_updates_1__din),
    .if_full_n(num_updates_1__full_n),
    .if_write(num_updates_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(49),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  num_updates_2
  (
    .clk(ap_clk),
    .reset(num_updates_2__rst__q2),
    .if_dout(num_updates_2__dout),
    .if_empty_n(num_updates_2__empty_n),
    .if_read(num_updates_2__read),
    .if_read_ce(1'b1),
    .if_din(num_updates_2__din),
    .if_full_n(num_updates_2__full_n),
    .if_write(num_updates_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(49),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  num_updates_3
  (
    .clk(ap_clk),
    .reset(num_updates_3__rst__q2),
    .if_dout(num_updates_3__dout),
    .if_empty_n(num_updates_3__empty_n),
    .if_read(num_updates_3__read),
    .if_read_ce(1'b1),
    .if_din(num_updates_3__din),
    .if_full_n(num_updates_3__full_n),
    .if_write(num_updates_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(49),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  num_updates_4
  (
    .clk(ap_clk),
    .reset(num_updates_4__rst__q2),
    .if_dout(num_updates_4__dout),
    .if_empty_n(num_updates_4__empty_n),
    .if_read(num_updates_4__read),
    .if_read_ce(1'b1),
    .if_din(num_updates_4__din),
    .if_full_n(num_updates_4__full_n),
    .if_write(num_updates_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(49),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  num_updates_5
  (
    .clk(ap_clk),
    .reset(num_updates_5__rst__q2),
    .if_dout(num_updates_5__dout),
    .if_empty_n(num_updates_5__empty_n),
    .if_read(num_updates_5__read),
    .if_read_ce(1'b1),
    .if_din(num_updates_5__din),
    .if_full_n(num_updates_5__full_n),
    .if_write(num_updates_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(49),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  num_updates_6
  (
    .clk(ap_clk),
    .reset(num_updates_6__rst__q2),
    .if_dout(num_updates_6__dout),
    .if_empty_n(num_updates_6__empty_n),
    .if_read(num_updates_6__read),
    .if_read_ce(1'b1),
    .if_din(num_updates_6__din),
    .if_full_n(num_updates_6__full_n),
    .if_write(num_updates_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(49),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  num_updates_7
  (
    .clk(ap_clk),
    .reset(num_updates_7__rst__q2),
    .if_dout(num_updates_7__dout),
    .if_empty_n(num_updates_7__empty_n),
    .if_read(num_updates_7__read),
    .if_read_ce(1'b1),
    .if_din(num_updates_7__din),
    .if_full_n(num_updates_7__full_n),
    .if_write(num_updates_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  scatter_phase_vertex_req
  (
    .clk(ap_clk),
    .reset(scatter_phase_vertex_req__rst__q2),
    .if_dout(scatter_phase_vertex_req__dout),
    .if_empty_n(scatter_phase_vertex_req__empty_n),
    .if_read(scatter_phase_vertex_req__read),
    .if_read_ce(1'b1),
    .if_din(scatter_phase_vertex_req__din),
    .if_full_n(scatter_phase_vertex_req__full_n),
    .if_write(scatter_phase_vertex_req__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(211),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_req_0
  (
    .clk(ap_clk),
    .reset(task_req_0__rst__q2),
    .if_dout(task_req_0__dout),
    .if_empty_n(task_req_0__empty_n),
    .if_read(task_req_0__read),
    .if_read_ce(1'b1),
    .if_din(task_req_0__din),
    .if_full_n(task_req_0__full_n),
    .if_write(task_req_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(211),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_req_1
  (
    .clk(ap_clk),
    .reset(task_req_1__rst__q2),
    .if_dout(task_req_1__dout),
    .if_empty_n(task_req_1__empty_n),
    .if_read(task_req_1__read),
    .if_read_ce(1'b1),
    .if_din(task_req_1__din),
    .if_full_n(task_req_1__full_n),
    .if_write(task_req_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(211),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_req_2
  (
    .clk(ap_clk),
    .reset(task_req_2__rst__q2),
    .if_dout(task_req_2__dout),
    .if_empty_n(task_req_2__empty_n),
    .if_read(task_req_2__read),
    .if_read_ce(1'b1),
    .if_din(task_req_2__din),
    .if_full_n(task_req_2__full_n),
    .if_write(task_req_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(211),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_req_3
  (
    .clk(ap_clk),
    .reset(task_req_3__rst__q2),
    .if_dout(task_req_3__dout),
    .if_empty_n(task_req_3__empty_n),
    .if_read(task_req_3__read),
    .if_read_ce(1'b1),
    .if_din(task_req_3__din),
    .if_full_n(task_req_3__full_n),
    .if_write(task_req_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(211),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_req_4
  (
    .clk(ap_clk),
    .reset(task_req_4__rst__q2),
    .if_dout(task_req_4__dout),
    .if_empty_n(task_req_4__empty_n),
    .if_read(task_req_4__read),
    .if_read_ce(1'b1),
    .if_din(task_req_4__din),
    .if_full_n(task_req_4__full_n),
    .if_write(task_req_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(211),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_req_5
  (
    .clk(ap_clk),
    .reset(task_req_5__rst__q2),
    .if_dout(task_req_5__dout),
    .if_empty_n(task_req_5__empty_n),
    .if_read(task_req_5__read),
    .if_read_ce(1'b1),
    .if_din(task_req_5__din),
    .if_full_n(task_req_5__full_n),
    .if_write(task_req_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(211),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_req_6
  (
    .clk(ap_clk),
    .reset(task_req_6__rst__q2),
    .if_dout(task_req_6__dout),
    .if_empty_n(task_req_6__empty_n),
    .if_read(task_req_6__read),
    .if_read_ce(1'b1),
    .if_din(task_req_6__din),
    .if_full_n(task_req_6__full_n),
    .if_write(task_req_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(211),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_req_7
  (
    .clk(ap_clk),
    .reset(task_req_7__rst__q2),
    .if_dout(task_req_7__dout),
    .if_empty_n(task_req_7__empty_n),
    .if_read(task_req_7__read),
    .if_read_ce(1'b1),
    .if_din(task_req_7__din),
    .if_full_n(task_req_7__full_n),
    .if_write(task_req_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_resp_0
  (
    .clk(ap_clk),
    .reset(task_resp_0__rst__q2),
    .if_dout(task_resp_0__dout),
    .if_empty_n(task_resp_0__empty_n),
    .if_read(task_resp_0__read),
    .if_read_ce(1'b1),
    .if_din(task_resp_0__din),
    .if_full_n(task_resp_0__full_n),
    .if_write(task_resp_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_resp_1
  (
    .clk(ap_clk),
    .reset(task_resp_1__rst__q2),
    .if_dout(task_resp_1__dout),
    .if_empty_n(task_resp_1__empty_n),
    .if_read(task_resp_1__read),
    .if_read_ce(1'b1),
    .if_din(task_resp_1__din),
    .if_full_n(task_resp_1__full_n),
    .if_write(task_resp_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_resp_2
  (
    .clk(ap_clk),
    .reset(task_resp_2__rst__q2),
    .if_dout(task_resp_2__dout),
    .if_empty_n(task_resp_2__empty_n),
    .if_read(task_resp_2__read),
    .if_read_ce(1'b1),
    .if_din(task_resp_2__din),
    .if_full_n(task_resp_2__full_n),
    .if_write(task_resp_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_resp_3
  (
    .clk(ap_clk),
    .reset(task_resp_3__rst__q2),
    .if_dout(task_resp_3__dout),
    .if_empty_n(task_resp_3__empty_n),
    .if_read(task_resp_3__read),
    .if_read_ce(1'b1),
    .if_din(task_resp_3__din),
    .if_full_n(task_resp_3__full_n),
    .if_write(task_resp_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_resp_4
  (
    .clk(ap_clk),
    .reset(task_resp_4__rst__q2),
    .if_dout(task_resp_4__dout),
    .if_empty_n(task_resp_4__empty_n),
    .if_read(task_resp_4__read),
    .if_read_ce(1'b1),
    .if_din(task_resp_4__din),
    .if_full_n(task_resp_4__full_n),
    .if_write(task_resp_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_resp_5
  (
    .clk(ap_clk),
    .reset(task_resp_5__rst__q2),
    .if_dout(task_resp_5__dout),
    .if_empty_n(task_resp_5__empty_n),
    .if_read(task_resp_5__read),
    .if_read_ce(1'b1),
    .if_din(task_resp_5__din),
    .if_full_n(task_resp_5__full_n),
    .if_write(task_resp_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_resp_6
  (
    .clk(ap_clk),
    .reset(task_resp_6__rst__q2),
    .if_dout(task_resp_6__dout),
    .if_empty_n(task_resp_6__empty_n),
    .if_read(task_resp_6__read),
    .if_read_ce(1'b1),
    .if_din(task_resp_6__din),
    .if_full_n(task_resp_6__full_n),
    .if_write(task_resp_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  task_resp_7
  (
    .clk(ap_clk),
    .reset(task_resp_7__rst__q2),
    .if_dout(task_resp_7__dout),
    .if_empty_n(task_resp_7__empty_n),
    .if_read(task_resp_7__read),
    .if_read_ce(1'b1),
    .if_din(task_resp_7__din),
    .if_full_n(task_resp_7__full_n),
    .if_write(task_resp_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_config_0
  (
    .clk(ap_clk),
    .reset(update_config_0__rst__q2),
    .if_dout(update_config_0__dout),
    .if_empty_n(update_config_0__empty_n),
    .if_read(update_config_0__read),
    .if_read_ce(1'b1),
    .if_din(update_config_0__din),
    .if_full_n(update_config_0__full_n),
    .if_write(update_config_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_config_1
  (
    .clk(ap_clk),
    .reset(update_config_1__rst__q2),
    .if_dout(update_config_1__dout),
    .if_empty_n(update_config_1__empty_n),
    .if_read(update_config_1__read),
    .if_read_ce(1'b1),
    .if_din(update_config_1__din),
    .if_full_n(update_config_1__full_n),
    .if_write(update_config_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_config_2
  (
    .clk(ap_clk),
    .reset(update_config_2__rst__q2),
    .if_dout(update_config_2__dout),
    .if_empty_n(update_config_2__empty_n),
    .if_read(update_config_2__read),
    .if_read_ce(1'b1),
    .if_din(update_config_2__din),
    .if_full_n(update_config_2__full_n),
    .if_write(update_config_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_config_3
  (
    .clk(ap_clk),
    .reset(update_config_3__rst__q2),
    .if_dout(update_config_3__dout),
    .if_empty_n(update_config_3__empty_n),
    .if_read(update_config_3__read),
    .if_read_ce(1'b1),
    .if_din(update_config_3__din),
    .if_full_n(update_config_3__full_n),
    .if_write(update_config_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_config_4
  (
    .clk(ap_clk),
    .reset(update_config_4__rst__q2),
    .if_dout(update_config_4__dout),
    .if_empty_n(update_config_4__empty_n),
    .if_read(update_config_4__read),
    .if_read_ce(1'b1),
    .if_din(update_config_4__din),
    .if_full_n(update_config_4__full_n),
    .if_write(update_config_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_config_5
  (
    .clk(ap_clk),
    .reset(update_config_5__rst__q2),
    .if_dout(update_config_5__dout),
    .if_empty_n(update_config_5__empty_n),
    .if_read(update_config_5__read),
    .if_read_ce(1'b1),
    .if_din(update_config_5__din),
    .if_full_n(update_config_5__full_n),
    .if_write(update_config_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_config_6
  (
    .clk(ap_clk),
    .reset(update_config_6__rst__q2),
    .if_dout(update_config_6__dout),
    .if_empty_n(update_config_6__empty_n),
    .if_read(update_config_6__read),
    .if_read_ce(1'b1),
    .if_din(update_config_6__din),
    .if_full_n(update_config_6__full_n),
    .if_write(update_config_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(33),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_config_7
  (
    .clk(ap_clk),
    .reset(update_config_7__rst__q2),
    .if_dout(update_config_7__dout),
    .if_empty_n(update_config_7__empty_n),
    .if_read(update_config_7__read),
    .if_read_ce(1'b1),
    .if_din(update_config_7__din),
    .if_full_n(update_config_7__full_n),
    .if_write(update_config_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_mm2pe_0
  (
    .clk(ap_clk),
    .reset(update_mm2pe_0__rst__q2),
    .if_dout(update_mm2pe_0__dout),
    .if_empty_n(update_mm2pe_0__empty_n),
    .if_read(update_mm2pe_0__read),
    .if_read_ce(1'b1),
    .if_din(update_mm2pe_0__din),
    .if_full_n(update_mm2pe_0__full_n),
    .if_write(update_mm2pe_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_mm2pe_1
  (
    .clk(ap_clk),
    .reset(update_mm2pe_1__rst__q2),
    .if_dout(update_mm2pe_1__dout),
    .if_empty_n(update_mm2pe_1__empty_n),
    .if_read(update_mm2pe_1__read),
    .if_read_ce(1'b1),
    .if_din(update_mm2pe_1__din),
    .if_full_n(update_mm2pe_1__full_n),
    .if_write(update_mm2pe_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_mm2pe_2
  (
    .clk(ap_clk),
    .reset(update_mm2pe_2__rst__q2),
    .if_dout(update_mm2pe_2__dout),
    .if_empty_n(update_mm2pe_2__empty_n),
    .if_read(update_mm2pe_2__read),
    .if_read_ce(1'b1),
    .if_din(update_mm2pe_2__din),
    .if_full_n(update_mm2pe_2__full_n),
    .if_write(update_mm2pe_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_mm2pe_3
  (
    .clk(ap_clk),
    .reset(update_mm2pe_3__rst__q2),
    .if_dout(update_mm2pe_3__dout),
    .if_empty_n(update_mm2pe_3__empty_n),
    .if_read(update_mm2pe_3__read),
    .if_read_ce(1'b1),
    .if_din(update_mm2pe_3__din),
    .if_full_n(update_mm2pe_3__full_n),
    .if_write(update_mm2pe_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_mm2pe_4
  (
    .clk(ap_clk),
    .reset(update_mm2pe_4__rst__q2),
    .if_dout(update_mm2pe_4__dout),
    .if_empty_n(update_mm2pe_4__empty_n),
    .if_read(update_mm2pe_4__read),
    .if_read_ce(1'b1),
    .if_din(update_mm2pe_4__din),
    .if_full_n(update_mm2pe_4__full_n),
    .if_write(update_mm2pe_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_mm2pe_5
  (
    .clk(ap_clk),
    .reset(update_mm2pe_5__rst__q2),
    .if_dout(update_mm2pe_5__dout),
    .if_empty_n(update_mm2pe_5__empty_n),
    .if_read(update_mm2pe_5__read),
    .if_read_ce(1'b1),
    .if_din(update_mm2pe_5__din),
    .if_full_n(update_mm2pe_5__full_n),
    .if_write(update_mm2pe_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_mm2pe_6
  (
    .clk(ap_clk),
    .reset(update_mm2pe_6__rst__q2),
    .if_dout(update_mm2pe_6__dout),
    .if_empty_n(update_mm2pe_6__empty_n),
    .if_read(update_mm2pe_6__read),
    .if_read_ce(1'b1),
    .if_din(update_mm2pe_6__din),
    .if_full_n(update_mm2pe_6__full_n),
    .if_write(update_mm2pe_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_mm2pe_7
  (
    .clk(ap_clk),
    .reset(update_mm2pe_7__rst__q2),
    .if_dout(update_mm2pe_7__dout),
    .if_empty_n(update_mm2pe_7__empty_n),
    .if_read(update_mm2pe_7__read),
    .if_read_ce(1'b1),
    .if_din(update_mm2pe_7__din),
    .if_full_n(update_mm2pe_7__full_n),
    .if_write(update_mm2pe_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(529),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_pe2mm_0
  (
    .clk(ap_clk),
    .reset(update_pe2mm_0__rst__q2),
    .if_dout(update_pe2mm_0__dout),
    .if_empty_n(update_pe2mm_0__empty_n),
    .if_read(update_pe2mm_0__read),
    .if_read_ce(1'b1),
    .if_din(update_pe2mm_0__din),
    .if_full_n(update_pe2mm_0__full_n),
    .if_write(update_pe2mm_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(529),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_pe2mm_1
  (
    .clk(ap_clk),
    .reset(update_pe2mm_1__rst__q2),
    .if_dout(update_pe2mm_1__dout),
    .if_empty_n(update_pe2mm_1__empty_n),
    .if_read(update_pe2mm_1__read),
    .if_read_ce(1'b1),
    .if_din(update_pe2mm_1__din),
    .if_full_n(update_pe2mm_1__full_n),
    .if_write(update_pe2mm_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(529),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_pe2mm_2
  (
    .clk(ap_clk),
    .reset(update_pe2mm_2__rst__q2),
    .if_dout(update_pe2mm_2__dout),
    .if_empty_n(update_pe2mm_2__empty_n),
    .if_read(update_pe2mm_2__read),
    .if_read_ce(1'b1),
    .if_din(update_pe2mm_2__din),
    .if_full_n(update_pe2mm_2__full_n),
    .if_write(update_pe2mm_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(529),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_pe2mm_3
  (
    .clk(ap_clk),
    .reset(update_pe2mm_3__rst__q2),
    .if_dout(update_pe2mm_3__dout),
    .if_empty_n(update_pe2mm_3__empty_n),
    .if_read(update_pe2mm_3__read),
    .if_read_ce(1'b1),
    .if_din(update_pe2mm_3__din),
    .if_full_n(update_pe2mm_3__full_n),
    .if_write(update_pe2mm_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(529),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_pe2mm_4
  (
    .clk(ap_clk),
    .reset(update_pe2mm_4__rst__q2),
    .if_dout(update_pe2mm_4__dout),
    .if_empty_n(update_pe2mm_4__empty_n),
    .if_read(update_pe2mm_4__read),
    .if_read_ce(1'b1),
    .if_din(update_pe2mm_4__din),
    .if_full_n(update_pe2mm_4__full_n),
    .if_write(update_pe2mm_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(529),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_pe2mm_5
  (
    .clk(ap_clk),
    .reset(update_pe2mm_5__rst__q2),
    .if_dout(update_pe2mm_5__dout),
    .if_empty_n(update_pe2mm_5__empty_n),
    .if_read(update_pe2mm_5__read),
    .if_read_ce(1'b1),
    .if_din(update_pe2mm_5__din),
    .if_full_n(update_pe2mm_5__full_n),
    .if_write(update_pe2mm_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(529),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_pe2mm_6
  (
    .clk(ap_clk),
    .reset(update_pe2mm_6__rst__q2),
    .if_dout(update_pe2mm_6__dout),
    .if_empty_n(update_pe2mm_6__empty_n),
    .if_read(update_pe2mm_6__read),
    .if_read_ce(1'b1),
    .if_din(update_pe2mm_6__din),
    .if_full_n(update_pe2mm_6__full_n),
    .if_write(update_pe2mm_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(529),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_pe2mm_7
  (
    .clk(ap_clk),
    .reset(update_pe2mm_7__rst__q2),
    .if_dout(update_pe2mm_7__dout),
    .if_empty_n(update_pe2mm_7__empty_n),
    .if_read(update_pe2mm_7__read),
    .if_read_ce(1'b1),
    .if_din(update_pe2mm_7__din),
    .if_full_n(update_pe2mm_7__full_n),
    .if_write(update_pe2mm_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_phase_0
  (
    .clk(ap_clk),
    .reset(update_phase_0__rst__q2),
    .if_dout(update_phase_0__dout),
    .if_empty_n(update_phase_0__empty_n),
    .if_read(update_phase_0__read),
    .if_read_ce(1'b1),
    .if_din(update_phase_0__din),
    .if_full_n(update_phase_0__full_n),
    .if_write(update_phase_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_phase_1
  (
    .clk(ap_clk),
    .reset(update_phase_1__rst__q2),
    .if_dout(update_phase_1__dout),
    .if_empty_n(update_phase_1__empty_n),
    .if_read(update_phase_1__read),
    .if_read_ce(1'b1),
    .if_din(update_phase_1__din),
    .if_full_n(update_phase_1__full_n),
    .if_write(update_phase_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_phase_2
  (
    .clk(ap_clk),
    .reset(update_phase_2__rst__q2),
    .if_dout(update_phase_2__dout),
    .if_empty_n(update_phase_2__empty_n),
    .if_read(update_phase_2__read),
    .if_read_ce(1'b1),
    .if_din(update_phase_2__din),
    .if_full_n(update_phase_2__full_n),
    .if_write(update_phase_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_phase_3
  (
    .clk(ap_clk),
    .reset(update_phase_3__rst__q2),
    .if_dout(update_phase_3__dout),
    .if_empty_n(update_phase_3__empty_n),
    .if_read(update_phase_3__read),
    .if_read_ce(1'b1),
    .if_din(update_phase_3__din),
    .if_full_n(update_phase_3__full_n),
    .if_write(update_phase_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_phase_4
  (
    .clk(ap_clk),
    .reset(update_phase_4__rst__q2),
    .if_dout(update_phase_4__dout),
    .if_empty_n(update_phase_4__empty_n),
    .if_read(update_phase_4__read),
    .if_read_ce(1'b1),
    .if_din(update_phase_4__din),
    .if_full_n(update_phase_4__full_n),
    .if_write(update_phase_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_phase_5
  (
    .clk(ap_clk),
    .reset(update_phase_5__rst__q2),
    .if_dout(update_phase_5__dout),
    .if_empty_n(update_phase_5__empty_n),
    .if_read(update_phase_5__read),
    .if_read_ce(1'b1),
    .if_din(update_phase_5__din),
    .if_full_n(update_phase_5__full_n),
    .if_write(update_phase_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_phase_6
  (
    .clk(ap_clk),
    .reset(update_phase_6__rst__q2),
    .if_dout(update_phase_6__dout),
    .if_empty_n(update_phase_6__empty_n),
    .if_read(update_phase_6__read),
    .if_read_ce(1'b1),
    .if_din(update_phase_6__din),
    .if_full_n(update_phase_6__full_n),
    .if_write(update_phase_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(2),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_phase_7
  (
    .clk(ap_clk),
    .reset(update_phase_7__rst__q2),
    .if_dout(update_phase_7__dout),
    .if_empty_n(update_phase_7__empty_n),
    .if_read(update_phase_7__read),
    .if_read_ce(1'b1),
    .if_din(update_phase_7__din),
    .if_full_n(update_phase_7__full_n),
    .if_write(update_phase_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_addr_0
  (
    .clk(ap_clk),
    .reset(update_read_addr_0__rst__q2),
    .if_dout(update_read_addr_0__dout),
    .if_empty_n(update_read_addr_0__empty_n),
    .if_read(update_read_addr_0__read),
    .if_read_ce(1'b1),
    .if_din(update_read_addr_0__din),
    .if_full_n(update_read_addr_0__full_n),
    .if_write(update_read_addr_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_addr_1
  (
    .clk(ap_clk),
    .reset(update_read_addr_1__rst__q2),
    .if_dout(update_read_addr_1__dout),
    .if_empty_n(update_read_addr_1__empty_n),
    .if_read(update_read_addr_1__read),
    .if_read_ce(1'b1),
    .if_din(update_read_addr_1__din),
    .if_full_n(update_read_addr_1__full_n),
    .if_write(update_read_addr_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_addr_2
  (
    .clk(ap_clk),
    .reset(update_read_addr_2__rst__q2),
    .if_dout(update_read_addr_2__dout),
    .if_empty_n(update_read_addr_2__empty_n),
    .if_read(update_read_addr_2__read),
    .if_read_ce(1'b1),
    .if_din(update_read_addr_2__din),
    .if_full_n(update_read_addr_2__full_n),
    .if_write(update_read_addr_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_addr_3
  (
    .clk(ap_clk),
    .reset(update_read_addr_3__rst__q2),
    .if_dout(update_read_addr_3__dout),
    .if_empty_n(update_read_addr_3__empty_n),
    .if_read(update_read_addr_3__read),
    .if_read_ce(1'b1),
    .if_din(update_read_addr_3__din),
    .if_full_n(update_read_addr_3__full_n),
    .if_write(update_read_addr_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_addr_4
  (
    .clk(ap_clk),
    .reset(update_read_addr_4__rst__q2),
    .if_dout(update_read_addr_4__dout),
    .if_empty_n(update_read_addr_4__empty_n),
    .if_read(update_read_addr_4__read),
    .if_read_ce(1'b1),
    .if_din(update_read_addr_4__din),
    .if_full_n(update_read_addr_4__full_n),
    .if_write(update_read_addr_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_addr_5
  (
    .clk(ap_clk),
    .reset(update_read_addr_5__rst__q2),
    .if_dout(update_read_addr_5__dout),
    .if_empty_n(update_read_addr_5__empty_n),
    .if_read(update_read_addr_5__read),
    .if_read_ce(1'b1),
    .if_din(update_read_addr_5__din),
    .if_full_n(update_read_addr_5__full_n),
    .if_write(update_read_addr_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_addr_6
  (
    .clk(ap_clk),
    .reset(update_read_addr_6__rst__q2),
    .if_dout(update_read_addr_6__dout),
    .if_empty_n(update_read_addr_6__empty_n),
    .if_read(update_read_addr_6__read),
    .if_read_ce(1'b1),
    .if_din(update_read_addr_6__din),
    .if_full_n(update_read_addr_6__full_n),
    .if_write(update_read_addr_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_addr_7
  (
    .clk(ap_clk),
    .reset(update_read_addr_7__rst__q2),
    .if_dout(update_read_addr_7__dout),
    .if_empty_n(update_read_addr_7__empty_n),
    .if_read(update_read_addr_7__read),
    .if_read_ce(1'b1),
    .if_din(update_read_addr_7__din),
    .if_full_n(update_read_addr_7__full_n),
    .if_write(update_read_addr_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_data_0
  (
    .clk(ap_clk),
    .reset(update_read_data_0__rst__q2),
    .if_dout(update_read_data_0__dout),
    .if_empty_n(update_read_data_0__empty_n),
    .if_read(update_read_data_0__read),
    .if_read_ce(1'b1),
    .if_din(update_read_data_0__din),
    .if_full_n(update_read_data_0__full_n),
    .if_write(update_read_data_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_data_1
  (
    .clk(ap_clk),
    .reset(update_read_data_1__rst__q2),
    .if_dout(update_read_data_1__dout),
    .if_empty_n(update_read_data_1__empty_n),
    .if_read(update_read_data_1__read),
    .if_read_ce(1'b1),
    .if_din(update_read_data_1__din),
    .if_full_n(update_read_data_1__full_n),
    .if_write(update_read_data_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_data_2
  (
    .clk(ap_clk),
    .reset(update_read_data_2__rst__q2),
    .if_dout(update_read_data_2__dout),
    .if_empty_n(update_read_data_2__empty_n),
    .if_read(update_read_data_2__read),
    .if_read_ce(1'b1),
    .if_din(update_read_data_2__din),
    .if_full_n(update_read_data_2__full_n),
    .if_write(update_read_data_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_data_3
  (
    .clk(ap_clk),
    .reset(update_read_data_3__rst__q2),
    .if_dout(update_read_data_3__dout),
    .if_empty_n(update_read_data_3__empty_n),
    .if_read(update_read_data_3__read),
    .if_read_ce(1'b1),
    .if_din(update_read_data_3__din),
    .if_full_n(update_read_data_3__full_n),
    .if_write(update_read_data_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_data_4
  (
    .clk(ap_clk),
    .reset(update_read_data_4__rst__q2),
    .if_dout(update_read_data_4__dout),
    .if_empty_n(update_read_data_4__empty_n),
    .if_read(update_read_data_4__read),
    .if_read_ce(1'b1),
    .if_din(update_read_data_4__din),
    .if_full_n(update_read_data_4__full_n),
    .if_write(update_read_data_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_data_5
  (
    .clk(ap_clk),
    .reset(update_read_data_5__rst__q2),
    .if_dout(update_read_data_5__dout),
    .if_empty_n(update_read_data_5__empty_n),
    .if_read(update_read_data_5__read),
    .if_read_ce(1'b1),
    .if_din(update_read_data_5__din),
    .if_full_n(update_read_data_5__full_n),
    .if_write(update_read_data_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_data_6
  (
    .clk(ap_clk),
    .reset(update_read_data_6__rst__q2),
    .if_dout(update_read_data_6__dout),
    .if_empty_n(update_read_data_6__empty_n),
    .if_read(update_read_data_6__read),
    .if_read_ce(1'b1),
    .if_din(update_read_data_6__din),
    .if_full_n(update_read_data_6__full_n),
    .if_write(update_read_data_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_read_data_7
  (
    .clk(ap_clk),
    .reset(update_read_data_7__rst__q2),
    .if_dout(update_read_data_7__dout),
    .if_empty_n(update_read_data_7__empty_n),
    .if_read(update_read_data_7__read),
    .if_read_ce(1'b1),
    .if_din(update_read_data_7__din),
    .if_full_n(update_read_data_7__full_n),
    .if_write(update_read_data_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(50),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_req_0
  (
    .clk(ap_clk),
    .reset(update_req_0__rst__q2),
    .if_dout(update_req_0__dout),
    .if_empty_n(update_req_0__empty_n),
    .if_read(update_req_0__read),
    .if_read_ce(1'b1),
    .if_din(update_req_0__din),
    .if_full_n(update_req_0__full_n),
    .if_write(update_req_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(50),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_req_1
  (
    .clk(ap_clk),
    .reset(update_req_1__rst__q2),
    .if_dout(update_req_1__dout),
    .if_empty_n(update_req_1__empty_n),
    .if_read(update_req_1__read),
    .if_read_ce(1'b1),
    .if_din(update_req_1__din),
    .if_full_n(update_req_1__full_n),
    .if_write(update_req_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(50),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_req_2
  (
    .clk(ap_clk),
    .reset(update_req_2__rst__q2),
    .if_dout(update_req_2__dout),
    .if_empty_n(update_req_2__empty_n),
    .if_read(update_req_2__read),
    .if_read_ce(1'b1),
    .if_din(update_req_2__din),
    .if_full_n(update_req_2__full_n),
    .if_write(update_req_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(50),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_req_3
  (
    .clk(ap_clk),
    .reset(update_req_3__rst__q2),
    .if_dout(update_req_3__dout),
    .if_empty_n(update_req_3__empty_n),
    .if_read(update_req_3__read),
    .if_read_ce(1'b1),
    .if_din(update_req_3__din),
    .if_full_n(update_req_3__full_n),
    .if_write(update_req_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(50),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_req_4
  (
    .clk(ap_clk),
    .reset(update_req_4__rst__q2),
    .if_dout(update_req_4__dout),
    .if_empty_n(update_req_4__empty_n),
    .if_read(update_req_4__read),
    .if_read_ce(1'b1),
    .if_din(update_req_4__din),
    .if_full_n(update_req_4__full_n),
    .if_write(update_req_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(50),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_req_5
  (
    .clk(ap_clk),
    .reset(update_req_5__rst__q2),
    .if_dout(update_req_5__dout),
    .if_empty_n(update_req_5__empty_n),
    .if_read(update_req_5__read),
    .if_read_ce(1'b1),
    .if_din(update_req_5__din),
    .if_full_n(update_req_5__full_n),
    .if_write(update_req_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(50),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_req_6
  (
    .clk(ap_clk),
    .reset(update_req_6__rst__q2),
    .if_dout(update_req_6__dout),
    .if_empty_n(update_req_6__empty_n),
    .if_read(update_req_6__read),
    .if_read_ce(1'b1),
    .if_din(update_req_6__din),
    .if_full_n(update_req_6__full_n),
    .if_write(update_req_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(50),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_req_7
  (
    .clk(ap_clk),
    .reset(update_req_7__rst__q2),
    .if_dout(update_req_7__dout),
    .if_empty_n(update_req_7__empty_n),
    .if_read(update_req_7__read),
    .if_read_ce(1'b1),
    .if_din(update_req_7__din),
    .if_full_n(update_req_7__full_n),
    .if_write(update_req_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_addr_0
  (
    .clk(ap_clk),
    .reset(update_write_addr_0__rst__q2),
    .if_dout(update_write_addr_0__dout),
    .if_empty_n(update_write_addr_0__empty_n),
    .if_read(update_write_addr_0__read),
    .if_read_ce(1'b1),
    .if_din(update_write_addr_0__din),
    .if_full_n(update_write_addr_0__full_n),
    .if_write(update_write_addr_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_addr_1
  (
    .clk(ap_clk),
    .reset(update_write_addr_1__rst__q2),
    .if_dout(update_write_addr_1__dout),
    .if_empty_n(update_write_addr_1__empty_n),
    .if_read(update_write_addr_1__read),
    .if_read_ce(1'b1),
    .if_din(update_write_addr_1__din),
    .if_full_n(update_write_addr_1__full_n),
    .if_write(update_write_addr_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_addr_2
  (
    .clk(ap_clk),
    .reset(update_write_addr_2__rst__q2),
    .if_dout(update_write_addr_2__dout),
    .if_empty_n(update_write_addr_2__empty_n),
    .if_read(update_write_addr_2__read),
    .if_read_ce(1'b1),
    .if_din(update_write_addr_2__din),
    .if_full_n(update_write_addr_2__full_n),
    .if_write(update_write_addr_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_addr_3
  (
    .clk(ap_clk),
    .reset(update_write_addr_3__rst__q2),
    .if_dout(update_write_addr_3__dout),
    .if_empty_n(update_write_addr_3__empty_n),
    .if_read(update_write_addr_3__read),
    .if_read_ce(1'b1),
    .if_din(update_write_addr_3__din),
    .if_full_n(update_write_addr_3__full_n),
    .if_write(update_write_addr_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_addr_4
  (
    .clk(ap_clk),
    .reset(update_write_addr_4__rst__q2),
    .if_dout(update_write_addr_4__dout),
    .if_empty_n(update_write_addr_4__empty_n),
    .if_read(update_write_addr_4__read),
    .if_read_ce(1'b1),
    .if_din(update_write_addr_4__din),
    .if_full_n(update_write_addr_4__full_n),
    .if_write(update_write_addr_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_addr_5
  (
    .clk(ap_clk),
    .reset(update_write_addr_5__rst__q2),
    .if_dout(update_write_addr_5__dout),
    .if_empty_n(update_write_addr_5__empty_n),
    .if_read(update_write_addr_5__read),
    .if_read_ce(1'b1),
    .if_din(update_write_addr_5__din),
    .if_full_n(update_write_addr_5__full_n),
    .if_write(update_write_addr_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_addr_6
  (
    .clk(ap_clk),
    .reset(update_write_addr_6__rst__q2),
    .if_dout(update_write_addr_6__dout),
    .if_empty_n(update_write_addr_6__empty_n),
    .if_read(update_write_addr_6__read),
    .if_read_ce(1'b1),
    .if_din(update_write_addr_6__din),
    .if_full_n(update_write_addr_6__full_n),
    .if_write(update_write_addr_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_addr_7
  (
    .clk(ap_clk),
    .reset(update_write_addr_7__rst__q2),
    .if_dout(update_write_addr_7__dout),
    .if_empty_n(update_write_addr_7__empty_n),
    .if_read(update_write_addr_7__read),
    .if_read_ce(1'b1),
    .if_din(update_write_addr_7__din),
    .if_full_n(update_write_addr_7__full_n),
    .if_write(update_write_addr_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_data_0
  (
    .clk(ap_clk),
    .reset(update_write_data_0__rst__q2),
    .if_dout(update_write_data_0__dout),
    .if_empty_n(update_write_data_0__empty_n),
    .if_read(update_write_data_0__read),
    .if_read_ce(1'b1),
    .if_din(update_write_data_0__din),
    .if_full_n(update_write_data_0__full_n),
    .if_write(update_write_data_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_data_1
  (
    .clk(ap_clk),
    .reset(update_write_data_1__rst__q2),
    .if_dout(update_write_data_1__dout),
    .if_empty_n(update_write_data_1__empty_n),
    .if_read(update_write_data_1__read),
    .if_read_ce(1'b1),
    .if_din(update_write_data_1__din),
    .if_full_n(update_write_data_1__full_n),
    .if_write(update_write_data_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_data_2
  (
    .clk(ap_clk),
    .reset(update_write_data_2__rst__q2),
    .if_dout(update_write_data_2__dout),
    .if_empty_n(update_write_data_2__empty_n),
    .if_read(update_write_data_2__read),
    .if_read_ce(1'b1),
    .if_din(update_write_data_2__din),
    .if_full_n(update_write_data_2__full_n),
    .if_write(update_write_data_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_data_3
  (
    .clk(ap_clk),
    .reset(update_write_data_3__rst__q2),
    .if_dout(update_write_data_3__dout),
    .if_empty_n(update_write_data_3__empty_n),
    .if_read(update_write_data_3__read),
    .if_read_ce(1'b1),
    .if_din(update_write_data_3__din),
    .if_full_n(update_write_data_3__full_n),
    .if_write(update_write_data_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_data_4
  (
    .clk(ap_clk),
    .reset(update_write_data_4__rst__q2),
    .if_dout(update_write_data_4__dout),
    .if_empty_n(update_write_data_4__empty_n),
    .if_read(update_write_data_4__read),
    .if_read_ce(1'b1),
    .if_din(update_write_data_4__din),
    .if_full_n(update_write_data_4__full_n),
    .if_write(update_write_data_4__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_data_5
  (
    .clk(ap_clk),
    .reset(update_write_data_5__rst__q2),
    .if_dout(update_write_data_5__dout),
    .if_empty_n(update_write_data_5__empty_n),
    .if_read(update_write_data_5__read),
    .if_read_ce(1'b1),
    .if_din(update_write_data_5__din),
    .if_full_n(update_write_data_5__full_n),
    .if_write(update_write_data_5__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_data_6
  (
    .clk(ap_clk),
    .reset(update_write_data_6__rst__q2),
    .if_dout(update_write_data_6__dout),
    .if_empty_n(update_write_data_6__empty_n),
    .if_read(update_write_data_6__read),
    .if_read_ce(1'b1),
    .if_din(update_write_data_6__din),
    .if_full_n(update_write_data_6__full_n),
    .if_write(update_write_data_6__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  update_write_data_7
  (
    .clk(ap_clk),
    .reset(update_write_data_7__rst__q2),
    .if_dout(update_write_data_7__dout),
    .if_empty_n(update_write_data_7__empty_n),
    .if_read(update_write_data_7__read),
    .if_read_ce(1'b1),
    .if_din(update_write_data_7__din),
    .if_full_n(update_write_data_7__full_n),
    .if_write(update_write_data_7__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r0_0
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r0_0__rst__q2),
    .if_dout(vertex_mm2pe_r0_0__dout),
    .if_empty_n(vertex_mm2pe_r0_0__empty_n),
    .if_read(vertex_mm2pe_r0_0__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r0_0__din),
    .if_full_n(vertex_mm2pe_r0_0__full_n),
    .if_write(vertex_mm2pe_r0_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r0_1
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r0_1__rst__q2),
    .if_dout(vertex_mm2pe_r0_1__dout),
    .if_empty_n(vertex_mm2pe_r0_1__empty_n),
    .if_read(vertex_mm2pe_r0_1__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r0_1__din),
    .if_full_n(vertex_mm2pe_r0_1__full_n),
    .if_write(vertex_mm2pe_r0_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r1_0
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r1_0__rst__q2),
    .if_dout(vertex_mm2pe_r1_0__dout),
    .if_empty_n(vertex_mm2pe_r1_0__empty_n),
    .if_read(vertex_mm2pe_r1_0__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r1_0__din),
    .if_full_n(vertex_mm2pe_r1_0__full_n),
    .if_write(vertex_mm2pe_r1_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r1_1
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r1_1__rst__q2),
    .if_dout(vertex_mm2pe_r1_1__dout),
    .if_empty_n(vertex_mm2pe_r1_1__empty_n),
    .if_read(vertex_mm2pe_r1_1__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r1_1__din),
    .if_full_n(vertex_mm2pe_r1_1__full_n),
    .if_write(vertex_mm2pe_r1_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r1_2
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r1_2__rst__q2),
    .if_dout(vertex_mm2pe_r1_2__dout),
    .if_empty_n(vertex_mm2pe_r1_2__empty_n),
    .if_read(vertex_mm2pe_r1_2__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r1_2__din),
    .if_full_n(vertex_mm2pe_r1_2__full_n),
    .if_write(vertex_mm2pe_r1_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r1_3
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r1_3__rst__q2),
    .if_dout(vertex_mm2pe_r1_3__dout),
    .if_empty_n(vertex_mm2pe_r1_3__empty_n),
    .if_read(vertex_mm2pe_r1_3__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r1_3__din),
    .if_full_n(vertex_mm2pe_r1_3__full_n),
    .if_write(vertex_mm2pe_r1_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r2_0
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r2_0__rst__q2),
    .if_dout(vertex_mm2pe_r2_0__dout),
    .if_empty_n(vertex_mm2pe_r2_0__empty_n),
    .if_read(vertex_mm2pe_r2_0__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r2_0__din),
    .if_full_n(vertex_mm2pe_r2_0__full_n),
    .if_write(vertex_mm2pe_r2_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r2_1
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r2_1__rst__q2),
    .if_dout(vertex_mm2pe_r2_1__dout),
    .if_empty_n(vertex_mm2pe_r2_1__empty_n),
    .if_read(vertex_mm2pe_r2_1__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r2_1__din),
    .if_full_n(vertex_mm2pe_r2_1__full_n),
    .if_write(vertex_mm2pe_r2_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r2_2
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r2_2__rst__q2),
    .if_dout(vertex_mm2pe_r2_2__dout),
    .if_empty_n(vertex_mm2pe_r2_2__empty_n),
    .if_read(vertex_mm2pe_r2_2__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r2_2__din),
    .if_full_n(vertex_mm2pe_r2_2__full_n),
    .if_write(vertex_mm2pe_r2_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_mm2pe_r2_3
  (
    .clk(ap_clk),
    .reset(vertex_mm2pe_r2_3__rst__q2),
    .if_dout(vertex_mm2pe_r2_3__dout),
    .if_empty_n(vertex_mm2pe_r2_3__empty_n),
    .if_read(vertex_mm2pe_r2_3__read),
    .if_read_ce(1'b1),
    .if_din(vertex_mm2pe_r2_3__din),
    .if_full_n(vertex_mm2pe_r2_3__full_n),
    .if_write(vertex_mm2pe_r2_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r0_0
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r0_0__rst__q2),
    .if_dout(vertex_pe2mm_r0_0__dout),
    .if_empty_n(vertex_pe2mm_r0_0__empty_n),
    .if_read(vertex_pe2mm_r0_0__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r0_0__din),
    .if_full_n(vertex_pe2mm_r0_0__full_n),
    .if_write(vertex_pe2mm_r0_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r0_1
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r0_1__rst__q2),
    .if_dout(vertex_pe2mm_r0_1__dout),
    .if_empty_n(vertex_pe2mm_r0_1__empty_n),
    .if_read(vertex_pe2mm_r0_1__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r0_1__din),
    .if_full_n(vertex_pe2mm_r0_1__full_n),
    .if_write(vertex_pe2mm_r0_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r1_0
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r1_0__rst__q2),
    .if_dout(vertex_pe2mm_r1_0__dout),
    .if_empty_n(vertex_pe2mm_r1_0__empty_n),
    .if_read(vertex_pe2mm_r1_0__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r1_0__din),
    .if_full_n(vertex_pe2mm_r1_0__full_n),
    .if_write(vertex_pe2mm_r1_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r1_1
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r1_1__rst__q2),
    .if_dout(vertex_pe2mm_r1_1__dout),
    .if_empty_n(vertex_pe2mm_r1_1__empty_n),
    .if_read(vertex_pe2mm_r1_1__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r1_1__din),
    .if_full_n(vertex_pe2mm_r1_1__full_n),
    .if_write(vertex_pe2mm_r1_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r1_2
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r1_2__rst__q2),
    .if_dout(vertex_pe2mm_r1_2__dout),
    .if_empty_n(vertex_pe2mm_r1_2__empty_n),
    .if_read(vertex_pe2mm_r1_2__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r1_2__din),
    .if_full_n(vertex_pe2mm_r1_2__full_n),
    .if_write(vertex_pe2mm_r1_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r1_3
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r1_3__rst__q2),
    .if_dout(vertex_pe2mm_r1_3__dout),
    .if_empty_n(vertex_pe2mm_r1_3__empty_n),
    .if_read(vertex_pe2mm_r1_3__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r1_3__din),
    .if_full_n(vertex_pe2mm_r1_3__full_n),
    .if_write(vertex_pe2mm_r1_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r2_0
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r2_0__rst__q2),
    .if_dout(vertex_pe2mm_r2_0__dout),
    .if_empty_n(vertex_pe2mm_r2_0__empty_n),
    .if_read(vertex_pe2mm_r2_0__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r2_0__din),
    .if_full_n(vertex_pe2mm_r2_0__full_n),
    .if_write(vertex_pe2mm_r2_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r2_1
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r2_1__rst__q2),
    .if_dout(vertex_pe2mm_r2_1__dout),
    .if_empty_n(vertex_pe2mm_r2_1__empty_n),
    .if_read(vertex_pe2mm_r2_1__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r2_1__din),
    .if_full_n(vertex_pe2mm_r2_1__full_n),
    .if_write(vertex_pe2mm_r2_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r2_2
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r2_2__rst__q2),
    .if_dout(vertex_pe2mm_r2_2__dout),
    .if_empty_n(vertex_pe2mm_r2_2__empty_n),
    .if_read(vertex_pe2mm_r2_2__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r2_2__din),
    .if_full_n(vertex_pe2mm_r2_2__full_n),
    .if_write(vertex_pe2mm_r2_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(1025),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_pe2mm_r2_3
  (
    .clk(ap_clk),
    .reset(vertex_pe2mm_r2_3__rst__q2),
    .if_dout(vertex_pe2mm_r2_3__dout),
    .if_empty_n(vertex_pe2mm_r2_3__empty_n),
    .if_read(vertex_pe2mm_r2_3__read),
    .if_read_ce(1'b1),
    .if_din(vertex_pe2mm_r2_3__din),
    .if_full_n(vertex_pe2mm_r2_3__full_n),
    .if_write(vertex_pe2mm_r2_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r0_0
  (
    .clk(ap_clk),
    .reset(vertex_req_r0_0__rst__q2),
    .if_dout(vertex_req_r0_0__dout),
    .if_empty_n(vertex_req_r0_0__empty_n),
    .if_read(vertex_req_r0_0__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r0_0__din),
    .if_full_n(vertex_req_r0_0__full_n),
    .if_write(vertex_req_r0_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r0_1
  (
    .clk(ap_clk),
    .reset(vertex_req_r0_1__rst__q2),
    .if_dout(vertex_req_r0_1__dout),
    .if_empty_n(vertex_req_r0_1__empty_n),
    .if_read(vertex_req_r0_1__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r0_1__din),
    .if_full_n(vertex_req_r0_1__full_n),
    .if_write(vertex_req_r0_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r1_0
  (
    .clk(ap_clk),
    .reset(vertex_req_r1_0__rst__q2),
    .if_dout(vertex_req_r1_0__dout),
    .if_empty_n(vertex_req_r1_0__empty_n),
    .if_read(vertex_req_r1_0__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r1_0__din),
    .if_full_n(vertex_req_r1_0__full_n),
    .if_write(vertex_req_r1_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r1_1
  (
    .clk(ap_clk),
    .reset(vertex_req_r1_1__rst__q2),
    .if_dout(vertex_req_r1_1__dout),
    .if_empty_n(vertex_req_r1_1__empty_n),
    .if_read(vertex_req_r1_1__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r1_1__din),
    .if_full_n(vertex_req_r1_1__full_n),
    .if_write(vertex_req_r1_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r1_2
  (
    .clk(ap_clk),
    .reset(vertex_req_r1_2__rst__q2),
    .if_dout(vertex_req_r1_2__dout),
    .if_empty_n(vertex_req_r1_2__empty_n),
    .if_read(vertex_req_r1_2__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r1_2__din),
    .if_full_n(vertex_req_r1_2__full_n),
    .if_write(vertex_req_r1_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r1_3
  (
    .clk(ap_clk),
    .reset(vertex_req_r1_3__rst__q2),
    .if_dout(vertex_req_r1_3__dout),
    .if_empty_n(vertex_req_r1_3__empty_n),
    .if_read(vertex_req_r1_3__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r1_3__din),
    .if_full_n(vertex_req_r1_3__full_n),
    .if_write(vertex_req_r1_3__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r2_0
  (
    .clk(ap_clk),
    .reset(vertex_req_r2_0__rst__q2),
    .if_dout(vertex_req_r2_0__dout),
    .if_empty_n(vertex_req_r2_0__empty_n),
    .if_read(vertex_req_r2_0__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r2_0__din),
    .if_full_n(vertex_req_r2_0__full_n),
    .if_write(vertex_req_r2_0__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r2_1
  (
    .clk(ap_clk),
    .reset(vertex_req_r2_1__rst__q2),
    .if_dout(vertex_req_r2_1__dout),
    .if_empty_n(vertex_req_r2_1__empty_n),
    .if_read(vertex_req_r2_1__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r2_1__din),
    .if_full_n(vertex_req_r2_1__full_n),
    .if_write(vertex_req_r2_1__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r2_2
  (
    .clk(ap_clk),
    .reset(vertex_req_r2_2__rst__q2),
    .if_dout(vertex_req_r2_2__dout),
    .if_empty_n(vertex_req_r2_2__empty_n),
    .if_read(vertex_req_r2_2__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r2_2__din),
    .if_full_n(vertex_req_r2_2__full_n),
    .if_write(vertex_req_r2_2__write),
    .if_write_ce(1'b1)
  );


  fifo
  #(
    .DATA_WIDTH(65),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  vertex_req_r2_3
  (
    .clk(ap_clk),
    .reset(vertex_req_r2_3__rst__q2),
    .if_dout(vertex_req_r2_3__dout),
    .if_empty_n(vertex_req_r2_3__empty_n),
    .if_read(vertex_req_r2_3__read),
    .if_read_ce(1'b1),
    .if_din(vertex_req_r2_3__din),
    .if_full_n(vertex_req_r2_3__full_n),
    .if_write(vertex_req_r2_3__write),
    .if_write_ce(1'b1)
  );


  Control_Control
  Control_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(Control_0__ap_rst_n__q2),
    .ap_start(Control_0__ap_start),
    .ap_done(Control_0__ap_done),
    .ap_idle(Control_0__ap_idle),
    .ap_ready(Control_0__ap_ready),
    .m_axi_metadata_ARADDR(m_axi_metadata_ARADDR),
    .m_axi_metadata_ARBURST(m_axi_metadata_ARBURST),
    .m_axi_metadata_ARCACHE(m_axi_metadata_ARCACHE),
    .m_axi_metadata_ARID(m_axi_metadata_ARID),
    .m_axi_metadata_ARLEN(m_axi_metadata_ARLEN),
    .m_axi_metadata_ARLOCK(m_axi_metadata_ARLOCK),
    .m_axi_metadata_ARPROT(m_axi_metadata_ARPROT),
    .m_axi_metadata_ARQOS(m_axi_metadata_ARQOS),
    .m_axi_metadata_ARREADY(m_axi_metadata_ARREADY),
    .m_axi_metadata_ARREGION(m_axi_metadata_ARREGION),
    .m_axi_metadata_ARSIZE(m_axi_metadata_ARSIZE),
    .m_axi_metadata_ARUSER(m_axi_metadata_ARUSER),
    .m_axi_metadata_ARVALID(m_axi_metadata_ARVALID),
    .m_axi_metadata_AWADDR(m_axi_metadata_AWADDR),
    .m_axi_metadata_AWBURST(m_axi_metadata_AWBURST),
    .m_axi_metadata_AWCACHE(m_axi_metadata_AWCACHE),
    .m_axi_metadata_AWID(m_axi_metadata_AWID),
    .m_axi_metadata_AWLEN(m_axi_metadata_AWLEN),
    .m_axi_metadata_AWLOCK(m_axi_metadata_AWLOCK),
    .m_axi_metadata_AWPROT(m_axi_metadata_AWPROT),
    .m_axi_metadata_AWQOS(m_axi_metadata_AWQOS),
    .m_axi_metadata_AWREADY(m_axi_metadata_AWREADY),
    .m_axi_metadata_AWREGION(m_axi_metadata_AWREGION),
    .m_axi_metadata_AWSIZE(m_axi_metadata_AWSIZE),
    .m_axi_metadata_AWUSER(m_axi_metadata_AWUSER),
    .m_axi_metadata_AWVALID(m_axi_metadata_AWVALID),
    .m_axi_metadata_BID(m_axi_metadata_BID),
    .m_axi_metadata_BREADY(m_axi_metadata_BREADY),
    .m_axi_metadata_BRESP(m_axi_metadata_BRESP),
    .m_axi_metadata_BUSER(m_axi_metadata_BUSER),
    .m_axi_metadata_BVALID(m_axi_metadata_BVALID),
    .m_axi_metadata_RDATA(m_axi_metadata_RDATA),
    .m_axi_metadata_RID(m_axi_metadata_RID),
    .m_axi_metadata_RLAST(m_axi_metadata_RLAST),
    .m_axi_metadata_RREADY(m_axi_metadata_RREADY),
    .m_axi_metadata_RRESP(m_axi_metadata_RRESP),
    .m_axi_metadata_RUSER(m_axi_metadata_RUSER),
    .m_axi_metadata_RVALID(m_axi_metadata_RVALID),
    .m_axi_metadata_WDATA(m_axi_metadata_WDATA),
    .m_axi_metadata_WID(m_axi_metadata_WID),
    .m_axi_metadata_WLAST(m_axi_metadata_WLAST),
    .m_axi_metadata_WREADY(m_axi_metadata_WREADY),
    .m_axi_metadata_WSTRB(m_axi_metadata_WSTRB),
    .m_axi_metadata_WUSER(m_axi_metadata_WUSER),
    .m_axi_metadata_WVALID(m_axi_metadata_WVALID),
    .metadata_offset(metadata__q2),
    .num_partitions(Control_0___num_partitions__q2),
    .num_updates_q_fifo_V_0_dout(num_updates_0__dout),
    .num_updates_q_fifo_V_0_empty_n(num_updates_0__empty_n),
    .num_updates_q_fifo_V_0_read(num_updates_0__read),
    .num_updates_q_peek_val_0(num_updates_0__dout),
    .num_updates_q_fifo_V_1_dout(num_updates_1__dout),
    .num_updates_q_fifo_V_1_empty_n(num_updates_1__empty_n),
    .num_updates_q_fifo_V_1_read(num_updates_1__read),
    .num_updates_q_peek_val_1(num_updates_1__dout),
    .num_updates_q_fifo_V_2_dout(num_updates_2__dout),
    .num_updates_q_fifo_V_2_empty_n(num_updates_2__empty_n),
    .num_updates_q_fifo_V_2_read(num_updates_2__read),
    .num_updates_q_peek_val_2(num_updates_2__dout),
    .num_updates_q_fifo_V_3_dout(num_updates_3__dout),
    .num_updates_q_fifo_V_3_empty_n(num_updates_3__empty_n),
    .num_updates_q_fifo_V_3_read(num_updates_3__read),
    .num_updates_q_peek_val_3(num_updates_3__dout),
    .num_updates_q_fifo_V_4_dout(num_updates_4__dout),
    .num_updates_q_fifo_V_4_empty_n(num_updates_4__empty_n),
    .num_updates_q_fifo_V_4_read(num_updates_4__read),
    .num_updates_q_peek_val_4(num_updates_4__dout),
    .num_updates_q_fifo_V_5_dout(num_updates_5__dout),
    .num_updates_q_fifo_V_5_empty_n(num_updates_5__empty_n),
    .num_updates_q_fifo_V_5_read(num_updates_5__read),
    .num_updates_q_peek_val_5(num_updates_5__dout),
    .num_updates_q_fifo_V_6_dout(num_updates_6__dout),
    .num_updates_q_fifo_V_6_empty_n(num_updates_6__empty_n),
    .num_updates_q_fifo_V_6_read(num_updates_6__read),
    .num_updates_q_peek_val_6(num_updates_6__dout),
    .num_updates_q_fifo_V_7_dout(num_updates_7__dout),
    .num_updates_q_fifo_V_7_empty_n(num_updates_7__empty_n),
    .num_updates_q_fifo_V_7_read(num_updates_7__read),
    .num_updates_q_peek_val_7(num_updates_7__dout),
    .vertex_req_q_fifo_V_din(scatter_phase_vertex_req__din),
    .vertex_req_q_fifo_V_full_n(scatter_phase_vertex_req__full_n),
    .vertex_req_q_fifo_V_write(scatter_phase_vertex_req__write),
    .task_req_q_fifo_V_0_din(task_req_0__din),
    .task_req_q_fifo_V_0_full_n(task_req_0__full_n),
    .task_req_q_fifo_V_0_write(task_req_0__write),
    .task_req_q_fifo_V_1_din(task_req_1__din),
    .task_req_q_fifo_V_1_full_n(task_req_1__full_n),
    .task_req_q_fifo_V_1_write(task_req_1__write),
    .task_req_q_fifo_V_2_din(task_req_2__din),
    .task_req_q_fifo_V_2_full_n(task_req_2__full_n),
    .task_req_q_fifo_V_2_write(task_req_2__write),
    .task_req_q_fifo_V_3_din(task_req_3__din),
    .task_req_q_fifo_V_3_full_n(task_req_3__full_n),
    .task_req_q_fifo_V_3_write(task_req_3__write),
    .task_req_q_fifo_V_4_din(task_req_4__din),
    .task_req_q_fifo_V_4_full_n(task_req_4__full_n),
    .task_req_q_fifo_V_4_write(task_req_4__write),
    .task_req_q_fifo_V_5_din(task_req_5__din),
    .task_req_q_fifo_V_5_full_n(task_req_5__full_n),
    .task_req_q_fifo_V_5_write(task_req_5__write),
    .task_req_q_fifo_V_6_din(task_req_6__din),
    .task_req_q_fifo_V_6_full_n(task_req_6__full_n),
    .task_req_q_fifo_V_6_write(task_req_6__write),
    .task_req_q_fifo_V_7_din(task_req_7__din),
    .task_req_q_fifo_V_7_full_n(task_req_7__full_n),
    .task_req_q_fifo_V_7_write(task_req_7__write),
    .task_resp_q_fifo_V_0_dout(task_resp_0__dout),
    .task_resp_q_fifo_V_0_empty_n(task_resp_0__empty_n),
    .task_resp_q_fifo_V_0_read(task_resp_0__read),
    .task_resp_q_peek_val_0(task_resp_0__dout),
    .task_resp_q_fifo_V_1_dout(task_resp_1__dout),
    .task_resp_q_fifo_V_1_empty_n(task_resp_1__empty_n),
    .task_resp_q_fifo_V_1_read(task_resp_1__read),
    .task_resp_q_peek_val_1(task_resp_1__dout),
    .task_resp_q_fifo_V_2_dout(task_resp_2__dout),
    .task_resp_q_fifo_V_2_empty_n(task_resp_2__empty_n),
    .task_resp_q_fifo_V_2_read(task_resp_2__read),
    .task_resp_q_peek_val_2(task_resp_2__dout),
    .task_resp_q_fifo_V_3_dout(task_resp_3__dout),
    .task_resp_q_fifo_V_3_empty_n(task_resp_3__empty_n),
    .task_resp_q_fifo_V_3_read(task_resp_3__read),
    .task_resp_q_peek_val_3(task_resp_3__dout),
    .task_resp_q_fifo_V_4_dout(task_resp_4__dout),
    .task_resp_q_fifo_V_4_empty_n(task_resp_4__empty_n),
    .task_resp_q_fifo_V_4_read(task_resp_4__read),
    .task_resp_q_peek_val_4(task_resp_4__dout),
    .task_resp_q_fifo_V_5_dout(task_resp_5__dout),
    .task_resp_q_fifo_V_5_empty_n(task_resp_5__empty_n),
    .task_resp_q_fifo_V_5_read(task_resp_5__read),
    .task_resp_q_peek_val_5(task_resp_5__dout),
    .task_resp_q_fifo_V_6_dout(task_resp_6__dout),
    .task_resp_q_fifo_V_6_empty_n(task_resp_6__empty_n),
    .task_resp_q_fifo_V_6_read(task_resp_6__read),
    .task_resp_q_peek_val_6(task_resp_6__dout),
    .task_resp_q_fifo_V_7_dout(task_resp_7__dout),
    .task_resp_q_fifo_V_7_empty_n(task_resp_7__empty_n),
    .task_resp_q_fifo_V_7_read(task_resp_7__read),
    .task_resp_q_peek_val_7(task_resp_7__dout),
    .update_config_q_fifo_V_0_din(update_config_0__din),
    .update_config_q_fifo_V_0_full_n(update_config_0__full_n),
    .update_config_q_fifo_V_0_write(update_config_0__write),
    .update_config_q_fifo_V_1_din(update_config_1__din),
    .update_config_q_fifo_V_1_full_n(update_config_1__full_n),
    .update_config_q_fifo_V_1_write(update_config_1__write),
    .update_config_q_fifo_V_2_din(update_config_2__din),
    .update_config_q_fifo_V_2_full_n(update_config_2__full_n),
    .update_config_q_fifo_V_2_write(update_config_2__write),
    .update_config_q_fifo_V_3_din(update_config_3__din),
    .update_config_q_fifo_V_3_full_n(update_config_3__full_n),
    .update_config_q_fifo_V_3_write(update_config_3__write),
    .update_config_q_fifo_V_4_din(update_config_4__din),
    .update_config_q_fifo_V_4_full_n(update_config_4__full_n),
    .update_config_q_fifo_V_4_write(update_config_4__write),
    .update_config_q_fifo_V_5_din(update_config_5__din),
    .update_config_q_fifo_V_5_full_n(update_config_5__full_n),
    .update_config_q_fifo_V_5_write(update_config_5__write),
    .update_config_q_fifo_V_6_din(update_config_6__din),
    .update_config_q_fifo_V_6_full_n(update_config_6__full_n),
    .update_config_q_fifo_V_6_write(update_config_6__write),
    .update_config_q_fifo_V_7_din(update_config_7__din),
    .update_config_q_fifo_V_7_full_n(update_config_7__full_n),
    .update_config_q_fifo_V_7_write(update_config_7__write),
    .update_phase_q_fifo_V_0_din(update_phase_0__din),
    .update_phase_q_fifo_V_0_full_n(update_phase_0__full_n),
    .update_phase_q_fifo_V_0_write(update_phase_0__write),
    .update_phase_q_fifo_V_1_din(update_phase_1__din),
    .update_phase_q_fifo_V_1_full_n(update_phase_1__full_n),
    .update_phase_q_fifo_V_1_write(update_phase_1__write),
    .update_phase_q_fifo_V_2_din(update_phase_2__din),
    .update_phase_q_fifo_V_2_full_n(update_phase_2__full_n),
    .update_phase_q_fifo_V_2_write(update_phase_2__write),
    .update_phase_q_fifo_V_3_din(update_phase_3__din),
    .update_phase_q_fifo_V_3_full_n(update_phase_3__full_n),
    .update_phase_q_fifo_V_3_write(update_phase_3__write),
    .update_phase_q_fifo_V_4_din(update_phase_4__din),
    .update_phase_q_fifo_V_4_full_n(update_phase_4__full_n),
    .update_phase_q_fifo_V_4_write(update_phase_4__write),
    .update_phase_q_fifo_V_5_din(update_phase_5__din),
    .update_phase_q_fifo_V_5_full_n(update_phase_5__full_n),
    .update_phase_q_fifo_V_5_write(update_phase_5__write),
    .update_phase_q_fifo_V_6_din(update_phase_6__din),
    .update_phase_q_fifo_V_6_full_n(update_phase_6__full_n),
    .update_phase_q_fifo_V_6_write(update_phase_6__write),
    .update_phase_q_fifo_V_7_din(update_phase_7__din),
    .update_phase_q_fifo_V_7_full_n(update_phase_7__full_n),
    .update_phase_q_fifo_V_7_write(update_phase_7__write)
  );


  EdgeMem_EdgeMem
  EdgeMem_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(EdgeMem_0__ap_rst_n__q2),
    .ap_start(EdgeMem_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .edge_req_q_fifo_V_dout(edge_req_0__dout),
    .edge_req_q_fifo_V_empty_n(edge_req_0__empty_n),
    .edge_req_q_fifo_V_read(edge_req_0__read),
    .edge_req_q_peek_val(edge_req_0__dout),
    .edge_resp_q_fifo_V_din(edge_resp_0__din),
    .edge_resp_q_fifo_V_full_n(edge_resp_0__full_n),
    .edge_resp_q_fifo_V_write(edge_resp_0__write),
    .edges_read_addr_V_din(edges_0_read_addr__din),
    .edges_read_addr_V_full_n(edges_0_read_addr__full_n),
    .edges_read_addr_V_write(edges_0_read_addr__write),
    .edges_read_data_V_data_V_dout(edges_0_read_data__dout),
    .edges_read_data_V_data_V_empty_n(edges_0_read_data__empty_n),
    .edges_read_data_V_data_V_read(edges_0_read_data__read)
  );


  EdgeMem_EdgeMem
  EdgeMem_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(EdgeMem_1__ap_rst_n__q2),
    .ap_start(EdgeMem_1__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .edge_req_q_fifo_V_dout(edge_req_1__dout),
    .edge_req_q_fifo_V_empty_n(edge_req_1__empty_n),
    .edge_req_q_fifo_V_read(edge_req_1__read),
    .edge_req_q_peek_val(edge_req_1__dout),
    .edge_resp_q_fifo_V_din(edge_resp_1__din),
    .edge_resp_q_fifo_V_full_n(edge_resp_1__full_n),
    .edge_resp_q_fifo_V_write(edge_resp_1__write),
    .edges_read_addr_V_din(edges_1_read_addr__din),
    .edges_read_addr_V_full_n(edges_1_read_addr__full_n),
    .edges_read_addr_V_write(edges_1_read_addr__write),
    .edges_read_data_V_data_V_dout(edges_1_read_data__dout),
    .edges_read_data_V_data_V_empty_n(edges_1_read_data__empty_n),
    .edges_read_data_V_data_V_read(edges_1_read_data__read)
  );


  EdgeMem_EdgeMem
  EdgeMem_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(EdgeMem_2__ap_rst_n__q2),
    .ap_start(EdgeMem_2__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .edge_req_q_fifo_V_dout(edge_req_2__dout),
    .edge_req_q_fifo_V_empty_n(edge_req_2__empty_n),
    .edge_req_q_fifo_V_read(edge_req_2__read),
    .edge_req_q_peek_val(edge_req_2__dout),
    .edge_resp_q_fifo_V_din(edge_resp_2__din),
    .edge_resp_q_fifo_V_full_n(edge_resp_2__full_n),
    .edge_resp_q_fifo_V_write(edge_resp_2__write),
    .edges_read_addr_V_din(edges_2_read_addr__din),
    .edges_read_addr_V_full_n(edges_2_read_addr__full_n),
    .edges_read_addr_V_write(edges_2_read_addr__write),
    .edges_read_data_V_data_V_dout(edges_2_read_data__dout),
    .edges_read_data_V_data_V_empty_n(edges_2_read_data__empty_n),
    .edges_read_data_V_data_V_read(edges_2_read_data__read)
  );


  EdgeMem_EdgeMem
  EdgeMem_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(EdgeMem_3__ap_rst_n__q2),
    .ap_start(EdgeMem_3__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .edge_req_q_fifo_V_dout(edge_req_3__dout),
    .edge_req_q_fifo_V_empty_n(edge_req_3__empty_n),
    .edge_req_q_fifo_V_read(edge_req_3__read),
    .edge_req_q_peek_val(edge_req_3__dout),
    .edge_resp_q_fifo_V_din(edge_resp_3__din),
    .edge_resp_q_fifo_V_full_n(edge_resp_3__full_n),
    .edge_resp_q_fifo_V_write(edge_resp_3__write),
    .edges_read_addr_V_din(edges_3_read_addr__din),
    .edges_read_addr_V_full_n(edges_3_read_addr__full_n),
    .edges_read_addr_V_write(edges_3_read_addr__write),
    .edges_read_data_V_data_V_dout(edges_3_read_data__dout),
    .edges_read_data_V_data_V_empty_n(edges_3_read_data__empty_n),
    .edges_read_data_V_data_V_read(edges_3_read_data__read)
  );


  EdgeMem_EdgeMem
  EdgeMem_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(EdgeMem_4__ap_rst_n__q2),
    .ap_start(EdgeMem_4__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .edge_req_q_fifo_V_dout(edge_req_4__dout),
    .edge_req_q_fifo_V_empty_n(edge_req_4__empty_n),
    .edge_req_q_fifo_V_read(edge_req_4__read),
    .edge_req_q_peek_val(edge_req_4__dout),
    .edge_resp_q_fifo_V_din(edge_resp_4__din),
    .edge_resp_q_fifo_V_full_n(edge_resp_4__full_n),
    .edge_resp_q_fifo_V_write(edge_resp_4__write),
    .edges_read_addr_V_din(edges_4_read_addr__din),
    .edges_read_addr_V_full_n(edges_4_read_addr__full_n),
    .edges_read_addr_V_write(edges_4_read_addr__write),
    .edges_read_data_V_data_V_dout(edges_4_read_data__dout),
    .edges_read_data_V_data_V_empty_n(edges_4_read_data__empty_n),
    .edges_read_data_V_data_V_read(edges_4_read_data__read)
  );


  EdgeMem_EdgeMem
  EdgeMem_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(EdgeMem_5__ap_rst_n__q2),
    .ap_start(EdgeMem_5__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .edge_req_q_fifo_V_dout(edge_req_5__dout),
    .edge_req_q_fifo_V_empty_n(edge_req_5__empty_n),
    .edge_req_q_fifo_V_read(edge_req_5__read),
    .edge_req_q_peek_val(edge_req_5__dout),
    .edge_resp_q_fifo_V_din(edge_resp_5__din),
    .edge_resp_q_fifo_V_full_n(edge_resp_5__full_n),
    .edge_resp_q_fifo_V_write(edge_resp_5__write),
    .edges_read_addr_V_din(edges_5_read_addr__din),
    .edges_read_addr_V_full_n(edges_5_read_addr__full_n),
    .edges_read_addr_V_write(edges_5_read_addr__write),
    .edges_read_data_V_data_V_dout(edges_5_read_data__dout),
    .edges_read_data_V_data_V_empty_n(edges_5_read_data__empty_n),
    .edges_read_data_V_data_V_read(edges_5_read_data__read)
  );


  EdgeMem_EdgeMem
  EdgeMem_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(EdgeMem_6__ap_rst_n__q2),
    .ap_start(EdgeMem_6__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .edge_req_q_fifo_V_dout(edge_req_6__dout),
    .edge_req_q_fifo_V_empty_n(edge_req_6__empty_n),
    .edge_req_q_fifo_V_read(edge_req_6__read),
    .edge_req_q_peek_val(edge_req_6__dout),
    .edge_resp_q_fifo_V_din(edge_resp_6__din),
    .edge_resp_q_fifo_V_full_n(edge_resp_6__full_n),
    .edge_resp_q_fifo_V_write(edge_resp_6__write),
    .edges_read_addr_V_din(edges_6_read_addr__din),
    .edges_read_addr_V_full_n(edges_6_read_addr__full_n),
    .edges_read_addr_V_write(edges_6_read_addr__write),
    .edges_read_data_V_data_V_dout(edges_6_read_data__dout),
    .edges_read_data_V_data_V_empty_n(edges_6_read_data__empty_n),
    .edges_read_data_V_data_V_read(edges_6_read_data__read)
  );


  EdgeMem_EdgeMem
  EdgeMem_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(EdgeMem_7__ap_rst_n__q2),
    .ap_start(EdgeMem_7__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .edge_req_q_fifo_V_dout(edge_req_7__dout),
    .edge_req_q_fifo_V_empty_n(edge_req_7__empty_n),
    .edge_req_q_fifo_V_read(edge_req_7__read),
    .edge_req_q_peek_val(edge_req_7__dout),
    .edge_resp_q_fifo_V_din(edge_resp_7__din),
    .edge_resp_q_fifo_V_full_n(edge_resp_7__full_n),
    .edge_resp_q_fifo_V_write(edge_resp_7__write),
    .edges_read_addr_V_din(edges_7_read_addr__din),
    .edges_read_addr_V_full_n(edges_7_read_addr__full_n),
    .edges_read_addr_V_write(edges_7_read_addr__write),
    .edges_read_data_V_data_V_dout(edges_7_read_data__dout),
    .edges_read_data_V_data_V_empty_n(edges_7_read_data__empty_n),
    .edges_read_data_V_data_V_read(edges_7_read_data__read)
  );


  ProcElem_ProcElem
  ProcElem_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ProcElem_0__ap_rst_n__q2),
    .ap_start(ProcElem_0__ap_start),
    .ap_done(ProcElem_0__ap_done),
    .ap_idle(ProcElem_0__ap_idle),
    .ap_ready(ProcElem_0__ap_ready),
    .edge_req_q_fifo_V_din(edge_req_0__din),
    .edge_req_q_fifo_V_full_n(edge_req_0__full_n),
    .edge_req_q_fifo_V_write(edge_req_0__write),
    .edge_resp_q_fifo_V_dout(edge_resp_0__dout),
    .edge_resp_q_fifo_V_empty_n(edge_resp_0__empty_n),
    .edge_resp_q_fifo_V_read(edge_resp_0__read),
    .edge_resp_q_peek_val(edge_resp_0__dout),
    .task_req_q_fifo_V_dout(task_req_0__dout),
    .task_req_q_fifo_V_empty_n(task_req_0__empty_n),
    .task_req_q_fifo_V_read(task_req_0__read),
    .task_req_q_peek_val(task_req_0__dout),
    .task_resp_q_fifo_V_din(task_resp_0__din),
    .task_resp_q_fifo_V_full_n(task_resp_0__full_n),
    .task_resp_q_fifo_V_write(task_resp_0__write),
    .update_in_q_fifo_V_dout(update_mm2pe_0__dout),
    .update_in_q_fifo_V_empty_n(update_mm2pe_0__empty_n),
    .update_in_q_fifo_V_read(update_mm2pe_0__read),
    .update_in_q_peek_val(update_mm2pe_0__dout),
    .update_out_q_fifo_V_din(update_pe2mm_0__din),
    .update_out_q_fifo_V_full_n(update_pe2mm_0__full_n),
    .update_out_q_fifo_V_write(update_pe2mm_0__write),
    .update_req_q_fifo_V_din(update_req_0__din),
    .update_req_q_fifo_V_full_n(update_req_0__full_n),
    .update_req_q_fifo_V_write(update_req_0__write),
    .vertex_in_q_fifo_V_dout(vertex_mm2pe_r0_0__dout),
    .vertex_in_q_fifo_V_empty_n(vertex_mm2pe_r0_0__empty_n),
    .vertex_in_q_fifo_V_read(vertex_mm2pe_r0_0__read),
    .vertex_in_q_peek_val(vertex_mm2pe_r0_0__dout),
    .vertex_out_q_fifo_V_din(vertex_pe2mm_r0_0__din),
    .vertex_out_q_fifo_V_full_n(vertex_pe2mm_r0_0__full_n),
    .vertex_out_q_fifo_V_write(vertex_pe2mm_r0_0__write),
    .vertex_req_q_fifo_V_din(vertex_req_r0_0__din),
    .vertex_req_q_fifo_V_full_n(vertex_req_r0_0__full_n),
    .vertex_req_q_fifo_V_write(vertex_req_r0_0__write)
  );


  ProcElem_ProcElem
  ProcElem_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ProcElem_1__ap_rst_n__q2),
    .ap_start(ProcElem_1__ap_start),
    .ap_done(ProcElem_1__ap_done),
    .ap_idle(ProcElem_1__ap_idle),
    .ap_ready(ProcElem_1__ap_ready),
    .edge_req_q_fifo_V_din(edge_req_1__din),
    .edge_req_q_fifo_V_full_n(edge_req_1__full_n),
    .edge_req_q_fifo_V_write(edge_req_1__write),
    .edge_resp_q_fifo_V_dout(edge_resp_1__dout),
    .edge_resp_q_fifo_V_empty_n(edge_resp_1__empty_n),
    .edge_resp_q_fifo_V_read(edge_resp_1__read),
    .edge_resp_q_peek_val(edge_resp_1__dout),
    .task_req_q_fifo_V_dout(task_req_1__dout),
    .task_req_q_fifo_V_empty_n(task_req_1__empty_n),
    .task_req_q_fifo_V_read(task_req_1__read),
    .task_req_q_peek_val(task_req_1__dout),
    .task_resp_q_fifo_V_din(task_resp_1__din),
    .task_resp_q_fifo_V_full_n(task_resp_1__full_n),
    .task_resp_q_fifo_V_write(task_resp_1__write),
    .update_in_q_fifo_V_dout(update_mm2pe_1__dout),
    .update_in_q_fifo_V_empty_n(update_mm2pe_1__empty_n),
    .update_in_q_fifo_V_read(update_mm2pe_1__read),
    .update_in_q_peek_val(update_mm2pe_1__dout),
    .update_out_q_fifo_V_din(update_pe2mm_1__din),
    .update_out_q_fifo_V_full_n(update_pe2mm_1__full_n),
    .update_out_q_fifo_V_write(update_pe2mm_1__write),
    .update_req_q_fifo_V_din(update_req_1__din),
    .update_req_q_fifo_V_full_n(update_req_1__full_n),
    .update_req_q_fifo_V_write(update_req_1__write),
    .vertex_in_q_fifo_V_dout(vertex_mm2pe_r1_0__dout),
    .vertex_in_q_fifo_V_empty_n(vertex_mm2pe_r1_0__empty_n),
    .vertex_in_q_fifo_V_read(vertex_mm2pe_r1_0__read),
    .vertex_in_q_peek_val(vertex_mm2pe_r1_0__dout),
    .vertex_out_q_fifo_V_din(vertex_pe2mm_r1_0__din),
    .vertex_out_q_fifo_V_full_n(vertex_pe2mm_r1_0__full_n),
    .vertex_out_q_fifo_V_write(vertex_pe2mm_r1_0__write),
    .vertex_req_q_fifo_V_din(vertex_req_r1_0__din),
    .vertex_req_q_fifo_V_full_n(vertex_req_r1_0__full_n),
    .vertex_req_q_fifo_V_write(vertex_req_r1_0__write)
  );


  ProcElem_ProcElem
  ProcElem_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ProcElem_2__ap_rst_n__q2),
    .ap_start(ProcElem_2__ap_start),
    .ap_done(ProcElem_2__ap_done),
    .ap_idle(ProcElem_2__ap_idle),
    .ap_ready(ProcElem_2__ap_ready),
    .edge_req_q_fifo_V_din(edge_req_2__din),
    .edge_req_q_fifo_V_full_n(edge_req_2__full_n),
    .edge_req_q_fifo_V_write(edge_req_2__write),
    .edge_resp_q_fifo_V_dout(edge_resp_2__dout),
    .edge_resp_q_fifo_V_empty_n(edge_resp_2__empty_n),
    .edge_resp_q_fifo_V_read(edge_resp_2__read),
    .edge_resp_q_peek_val(edge_resp_2__dout),
    .task_req_q_fifo_V_dout(task_req_2__dout),
    .task_req_q_fifo_V_empty_n(task_req_2__empty_n),
    .task_req_q_fifo_V_read(task_req_2__read),
    .task_req_q_peek_val(task_req_2__dout),
    .task_resp_q_fifo_V_din(task_resp_2__din),
    .task_resp_q_fifo_V_full_n(task_resp_2__full_n),
    .task_resp_q_fifo_V_write(task_resp_2__write),
    .update_in_q_fifo_V_dout(update_mm2pe_2__dout),
    .update_in_q_fifo_V_empty_n(update_mm2pe_2__empty_n),
    .update_in_q_fifo_V_read(update_mm2pe_2__read),
    .update_in_q_peek_val(update_mm2pe_2__dout),
    .update_out_q_fifo_V_din(update_pe2mm_2__din),
    .update_out_q_fifo_V_full_n(update_pe2mm_2__full_n),
    .update_out_q_fifo_V_write(update_pe2mm_2__write),
    .update_req_q_fifo_V_din(update_req_2__din),
    .update_req_q_fifo_V_full_n(update_req_2__full_n),
    .update_req_q_fifo_V_write(update_req_2__write),
    .vertex_in_q_fifo_V_dout(vertex_mm2pe_r1_1__dout),
    .vertex_in_q_fifo_V_empty_n(vertex_mm2pe_r1_1__empty_n),
    .vertex_in_q_fifo_V_read(vertex_mm2pe_r1_1__read),
    .vertex_in_q_peek_val(vertex_mm2pe_r1_1__dout),
    .vertex_out_q_fifo_V_din(vertex_pe2mm_r1_1__din),
    .vertex_out_q_fifo_V_full_n(vertex_pe2mm_r1_1__full_n),
    .vertex_out_q_fifo_V_write(vertex_pe2mm_r1_1__write),
    .vertex_req_q_fifo_V_din(vertex_req_r1_1__din),
    .vertex_req_q_fifo_V_full_n(vertex_req_r1_1__full_n),
    .vertex_req_q_fifo_V_write(vertex_req_r1_1__write)
  );


  ProcElem_ProcElem
  ProcElem_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ProcElem_3__ap_rst_n__q2),
    .ap_start(ProcElem_3__ap_start),
    .ap_done(ProcElem_3__ap_done),
    .ap_idle(ProcElem_3__ap_idle),
    .ap_ready(ProcElem_3__ap_ready),
    .edge_req_q_fifo_V_din(edge_req_3__din),
    .edge_req_q_fifo_V_full_n(edge_req_3__full_n),
    .edge_req_q_fifo_V_write(edge_req_3__write),
    .edge_resp_q_fifo_V_dout(edge_resp_3__dout),
    .edge_resp_q_fifo_V_empty_n(edge_resp_3__empty_n),
    .edge_resp_q_fifo_V_read(edge_resp_3__read),
    .edge_resp_q_peek_val(edge_resp_3__dout),
    .task_req_q_fifo_V_dout(task_req_3__dout),
    .task_req_q_fifo_V_empty_n(task_req_3__empty_n),
    .task_req_q_fifo_V_read(task_req_3__read),
    .task_req_q_peek_val(task_req_3__dout),
    .task_resp_q_fifo_V_din(task_resp_3__din),
    .task_resp_q_fifo_V_full_n(task_resp_3__full_n),
    .task_resp_q_fifo_V_write(task_resp_3__write),
    .update_in_q_fifo_V_dout(update_mm2pe_3__dout),
    .update_in_q_fifo_V_empty_n(update_mm2pe_3__empty_n),
    .update_in_q_fifo_V_read(update_mm2pe_3__read),
    .update_in_q_peek_val(update_mm2pe_3__dout),
    .update_out_q_fifo_V_din(update_pe2mm_3__din),
    .update_out_q_fifo_V_full_n(update_pe2mm_3__full_n),
    .update_out_q_fifo_V_write(update_pe2mm_3__write),
    .update_req_q_fifo_V_din(update_req_3__din),
    .update_req_q_fifo_V_full_n(update_req_3__full_n),
    .update_req_q_fifo_V_write(update_req_3__write),
    .vertex_in_q_fifo_V_dout(vertex_mm2pe_r1_2__dout),
    .vertex_in_q_fifo_V_empty_n(vertex_mm2pe_r1_2__empty_n),
    .vertex_in_q_fifo_V_read(vertex_mm2pe_r1_2__read),
    .vertex_in_q_peek_val(vertex_mm2pe_r1_2__dout),
    .vertex_out_q_fifo_V_din(vertex_pe2mm_r1_2__din),
    .vertex_out_q_fifo_V_full_n(vertex_pe2mm_r1_2__full_n),
    .vertex_out_q_fifo_V_write(vertex_pe2mm_r1_2__write),
    .vertex_req_q_fifo_V_din(vertex_req_r1_2__din),
    .vertex_req_q_fifo_V_full_n(vertex_req_r1_2__full_n),
    .vertex_req_q_fifo_V_write(vertex_req_r1_2__write)
  );


  ProcElem_ProcElem
  ProcElem_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ProcElem_4__ap_rst_n__q2),
    .ap_start(ProcElem_4__ap_start),
    .ap_done(ProcElem_4__ap_done),
    .ap_idle(ProcElem_4__ap_idle),
    .ap_ready(ProcElem_4__ap_ready),
    .edge_req_q_fifo_V_din(edge_req_4__din),
    .edge_req_q_fifo_V_full_n(edge_req_4__full_n),
    .edge_req_q_fifo_V_write(edge_req_4__write),
    .edge_resp_q_fifo_V_dout(edge_resp_4__dout),
    .edge_resp_q_fifo_V_empty_n(edge_resp_4__empty_n),
    .edge_resp_q_fifo_V_read(edge_resp_4__read),
    .edge_resp_q_peek_val(edge_resp_4__dout),
    .task_req_q_fifo_V_dout(task_req_4__dout),
    .task_req_q_fifo_V_empty_n(task_req_4__empty_n),
    .task_req_q_fifo_V_read(task_req_4__read),
    .task_req_q_peek_val(task_req_4__dout),
    .task_resp_q_fifo_V_din(task_resp_4__din),
    .task_resp_q_fifo_V_full_n(task_resp_4__full_n),
    .task_resp_q_fifo_V_write(task_resp_4__write),
    .update_in_q_fifo_V_dout(update_mm2pe_4__dout),
    .update_in_q_fifo_V_empty_n(update_mm2pe_4__empty_n),
    .update_in_q_fifo_V_read(update_mm2pe_4__read),
    .update_in_q_peek_val(update_mm2pe_4__dout),
    .update_out_q_fifo_V_din(update_pe2mm_4__din),
    .update_out_q_fifo_V_full_n(update_pe2mm_4__full_n),
    .update_out_q_fifo_V_write(update_pe2mm_4__write),
    .update_req_q_fifo_V_din(update_req_4__din),
    .update_req_q_fifo_V_full_n(update_req_4__full_n),
    .update_req_q_fifo_V_write(update_req_4__write),
    .vertex_in_q_fifo_V_dout(vertex_mm2pe_r2_0__dout),
    .vertex_in_q_fifo_V_empty_n(vertex_mm2pe_r2_0__empty_n),
    .vertex_in_q_fifo_V_read(vertex_mm2pe_r2_0__read),
    .vertex_in_q_peek_val(vertex_mm2pe_r2_0__dout),
    .vertex_out_q_fifo_V_din(vertex_pe2mm_r2_0__din),
    .vertex_out_q_fifo_V_full_n(vertex_pe2mm_r2_0__full_n),
    .vertex_out_q_fifo_V_write(vertex_pe2mm_r2_0__write),
    .vertex_req_q_fifo_V_din(vertex_req_r2_0__din),
    .vertex_req_q_fifo_V_full_n(vertex_req_r2_0__full_n),
    .vertex_req_q_fifo_V_write(vertex_req_r2_0__write)
  );


  ProcElem_ProcElem
  ProcElem_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ProcElem_5__ap_rst_n__q2),
    .ap_start(ProcElem_5__ap_start),
    .ap_done(ProcElem_5__ap_done),
    .ap_idle(ProcElem_5__ap_idle),
    .ap_ready(ProcElem_5__ap_ready),
    .edge_req_q_fifo_V_din(edge_req_5__din),
    .edge_req_q_fifo_V_full_n(edge_req_5__full_n),
    .edge_req_q_fifo_V_write(edge_req_5__write),
    .edge_resp_q_fifo_V_dout(edge_resp_5__dout),
    .edge_resp_q_fifo_V_empty_n(edge_resp_5__empty_n),
    .edge_resp_q_fifo_V_read(edge_resp_5__read),
    .edge_resp_q_peek_val(edge_resp_5__dout),
    .task_req_q_fifo_V_dout(task_req_5__dout),
    .task_req_q_fifo_V_empty_n(task_req_5__empty_n),
    .task_req_q_fifo_V_read(task_req_5__read),
    .task_req_q_peek_val(task_req_5__dout),
    .task_resp_q_fifo_V_din(task_resp_5__din),
    .task_resp_q_fifo_V_full_n(task_resp_5__full_n),
    .task_resp_q_fifo_V_write(task_resp_5__write),
    .update_in_q_fifo_V_dout(update_mm2pe_5__dout),
    .update_in_q_fifo_V_empty_n(update_mm2pe_5__empty_n),
    .update_in_q_fifo_V_read(update_mm2pe_5__read),
    .update_in_q_peek_val(update_mm2pe_5__dout),
    .update_out_q_fifo_V_din(update_pe2mm_5__din),
    .update_out_q_fifo_V_full_n(update_pe2mm_5__full_n),
    .update_out_q_fifo_V_write(update_pe2mm_5__write),
    .update_req_q_fifo_V_din(update_req_5__din),
    .update_req_q_fifo_V_full_n(update_req_5__full_n),
    .update_req_q_fifo_V_write(update_req_5__write),
    .vertex_in_q_fifo_V_dout(vertex_mm2pe_r2_1__dout),
    .vertex_in_q_fifo_V_empty_n(vertex_mm2pe_r2_1__empty_n),
    .vertex_in_q_fifo_V_read(vertex_mm2pe_r2_1__read),
    .vertex_in_q_peek_val(vertex_mm2pe_r2_1__dout),
    .vertex_out_q_fifo_V_din(vertex_pe2mm_r2_1__din),
    .vertex_out_q_fifo_V_full_n(vertex_pe2mm_r2_1__full_n),
    .vertex_out_q_fifo_V_write(vertex_pe2mm_r2_1__write),
    .vertex_req_q_fifo_V_din(vertex_req_r2_1__din),
    .vertex_req_q_fifo_V_full_n(vertex_req_r2_1__full_n),
    .vertex_req_q_fifo_V_write(vertex_req_r2_1__write)
  );


  ProcElem_ProcElem
  ProcElem_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ProcElem_6__ap_rst_n__q2),
    .ap_start(ProcElem_6__ap_start),
    .ap_done(ProcElem_6__ap_done),
    .ap_idle(ProcElem_6__ap_idle),
    .ap_ready(ProcElem_6__ap_ready),
    .edge_req_q_fifo_V_din(edge_req_6__din),
    .edge_req_q_fifo_V_full_n(edge_req_6__full_n),
    .edge_req_q_fifo_V_write(edge_req_6__write),
    .edge_resp_q_fifo_V_dout(edge_resp_6__dout),
    .edge_resp_q_fifo_V_empty_n(edge_resp_6__empty_n),
    .edge_resp_q_fifo_V_read(edge_resp_6__read),
    .edge_resp_q_peek_val(edge_resp_6__dout),
    .task_req_q_fifo_V_dout(task_req_6__dout),
    .task_req_q_fifo_V_empty_n(task_req_6__empty_n),
    .task_req_q_fifo_V_read(task_req_6__read),
    .task_req_q_peek_val(task_req_6__dout),
    .task_resp_q_fifo_V_din(task_resp_6__din),
    .task_resp_q_fifo_V_full_n(task_resp_6__full_n),
    .task_resp_q_fifo_V_write(task_resp_6__write),
    .update_in_q_fifo_V_dout(update_mm2pe_6__dout),
    .update_in_q_fifo_V_empty_n(update_mm2pe_6__empty_n),
    .update_in_q_fifo_V_read(update_mm2pe_6__read),
    .update_in_q_peek_val(update_mm2pe_6__dout),
    .update_out_q_fifo_V_din(update_pe2mm_6__din),
    .update_out_q_fifo_V_full_n(update_pe2mm_6__full_n),
    .update_out_q_fifo_V_write(update_pe2mm_6__write),
    .update_req_q_fifo_V_din(update_req_6__din),
    .update_req_q_fifo_V_full_n(update_req_6__full_n),
    .update_req_q_fifo_V_write(update_req_6__write),
    .vertex_in_q_fifo_V_dout(vertex_mm2pe_r2_2__dout),
    .vertex_in_q_fifo_V_empty_n(vertex_mm2pe_r2_2__empty_n),
    .vertex_in_q_fifo_V_read(vertex_mm2pe_r2_2__read),
    .vertex_in_q_peek_val(vertex_mm2pe_r2_2__dout),
    .vertex_out_q_fifo_V_din(vertex_pe2mm_r2_2__din),
    .vertex_out_q_fifo_V_full_n(vertex_pe2mm_r2_2__full_n),
    .vertex_out_q_fifo_V_write(vertex_pe2mm_r2_2__write),
    .vertex_req_q_fifo_V_din(vertex_req_r2_2__din),
    .vertex_req_q_fifo_V_full_n(vertex_req_r2_2__full_n),
    .vertex_req_q_fifo_V_write(vertex_req_r2_2__write)
  );


  ProcElem_ProcElem
  ProcElem_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ProcElem_7__ap_rst_n__q2),
    .ap_start(ProcElem_7__ap_start),
    .ap_done(ProcElem_7__ap_done),
    .ap_idle(ProcElem_7__ap_idle),
    .ap_ready(ProcElem_7__ap_ready),
    .edge_req_q_fifo_V_din(edge_req_7__din),
    .edge_req_q_fifo_V_full_n(edge_req_7__full_n),
    .edge_req_q_fifo_V_write(edge_req_7__write),
    .edge_resp_q_fifo_V_dout(edge_resp_7__dout),
    .edge_resp_q_fifo_V_empty_n(edge_resp_7__empty_n),
    .edge_resp_q_fifo_V_read(edge_resp_7__read),
    .edge_resp_q_peek_val(edge_resp_7__dout),
    .task_req_q_fifo_V_dout(task_req_7__dout),
    .task_req_q_fifo_V_empty_n(task_req_7__empty_n),
    .task_req_q_fifo_V_read(task_req_7__read),
    .task_req_q_peek_val(task_req_7__dout),
    .task_resp_q_fifo_V_din(task_resp_7__din),
    .task_resp_q_fifo_V_full_n(task_resp_7__full_n),
    .task_resp_q_fifo_V_write(task_resp_7__write),
    .update_in_q_fifo_V_dout(update_mm2pe_7__dout),
    .update_in_q_fifo_V_empty_n(update_mm2pe_7__empty_n),
    .update_in_q_fifo_V_read(update_mm2pe_7__read),
    .update_in_q_peek_val(update_mm2pe_7__dout),
    .update_out_q_fifo_V_din(update_pe2mm_7__din),
    .update_out_q_fifo_V_full_n(update_pe2mm_7__full_n),
    .update_out_q_fifo_V_write(update_pe2mm_7__write),
    .update_req_q_fifo_V_din(update_req_7__din),
    .update_req_q_fifo_V_full_n(update_req_7__full_n),
    .update_req_q_fifo_V_write(update_req_7__write),
    .vertex_in_q_fifo_V_dout(vertex_mm2pe_r2_3__dout),
    .vertex_in_q_fifo_V_empty_n(vertex_mm2pe_r2_3__empty_n),
    .vertex_in_q_fifo_V_read(vertex_mm2pe_r2_3__read),
    .vertex_in_q_peek_val(vertex_mm2pe_r2_3__dout),
    .vertex_out_q_fifo_V_din(vertex_pe2mm_r2_3__din),
    .vertex_out_q_fifo_V_full_n(vertex_pe2mm_r2_3__full_n),
    .vertex_out_q_fifo_V_write(vertex_pe2mm_r2_3__write),
    .vertex_req_q_fifo_V_din(vertex_req_r2_3__din),
    .vertex_req_q_fifo_V_full_n(vertex_req_r2_3__full_n),
    .vertex_req_q_fifo_V_write(vertex_req_r2_3__write)
  );


  UpdateHandler_UpdateHandler
  UpdateHandler_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateHandler_0__ap_rst_n__q2),
    .ap_start(UpdateHandler_0__ap_start),
    .ap_done(UpdateHandler_0__ap_done),
    .ap_idle(UpdateHandler_0__ap_idle),
    .ap_ready(UpdateHandler_0__ap_ready),
    .num_partitions(UpdateHandler_0___num_partitions__q2),
    .num_updates_out_q_fifo_V_din(num_updates_0__din),
    .num_updates_out_q_fifo_V_full_n(num_updates_0__full_n),
    .num_updates_out_q_fifo_V_write(num_updates_0__write),
    .update_config_q_fifo_V_dout(update_config_0__dout),
    .update_config_q_fifo_V_empty_n(update_config_0__empty_n),
    .update_config_q_fifo_V_read(update_config_0__read),
    .update_config_q_peek_val(update_config_0__dout),
    .update_out_q_fifo_V_din(update_mm2pe_0__din),
    .update_out_q_fifo_V_full_n(update_mm2pe_0__full_n),
    .update_out_q_fifo_V_write(update_mm2pe_0__write),
    .update_in_q_fifo_V_dout(update_pe2mm_0__dout),
    .update_in_q_fifo_V_empty_n(update_pe2mm_0__empty_n),
    .update_in_q_fifo_V_read(update_pe2mm_0__read),
    .update_in_q_peek_val(update_pe2mm_0__dout),
    .update_phase_q_fifo_V_dout(update_phase_0__dout),
    .update_phase_q_fifo_V_empty_n(update_phase_0__empty_n),
    .update_phase_q_fifo_V_read(update_phase_0__read),
    .update_phase_q_peek_val(update_phase_0__dout),
    .updates_read_addr_q_fifo_V_din(update_read_addr_0__din),
    .updates_read_addr_q_fifo_V_full_n(update_read_addr_0__full_n),
    .updates_read_addr_q_fifo_V_write(update_read_addr_0__write),
    .updates_read_data_q_fifo_V_dout(update_read_data_0__dout),
    .updates_read_data_q_fifo_V_empty_n(update_read_data_0__empty_n),
    .updates_read_data_q_fifo_V_read(update_read_data_0__read),
    .updates_read_data_q_peek_val(update_read_data_0__dout),
    .update_req_q_fifo_V_dout(update_req_0__dout),
    .update_req_q_fifo_V_empty_n(update_req_0__empty_n),
    .update_req_q_fifo_V_read(update_req_0__read),
    .update_req_q_peek_val(update_req_0__dout),
    .updates_write_addr_q_fifo_V_din(update_write_addr_0__din),
    .updates_write_addr_q_fifo_V_full_n(update_write_addr_0__full_n),
    .updates_write_addr_q_fifo_V_write(update_write_addr_0__write),
    .updates_write_data_q_fifo_V_din(update_write_data_0__din),
    .updates_write_data_q_fifo_V_full_n(update_write_data_0__full_n),
    .updates_write_data_q_fifo_V_write(update_write_data_0__write)
  );


  UpdateHandler_UpdateHandler
  UpdateHandler_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateHandler_1__ap_rst_n__q2),
    .ap_start(UpdateHandler_1__ap_start),
    .ap_done(UpdateHandler_1__ap_done),
    .ap_idle(UpdateHandler_1__ap_idle),
    .ap_ready(UpdateHandler_1__ap_ready),
    .num_partitions(UpdateHandler_1___num_partitions__q2),
    .num_updates_out_q_fifo_V_din(num_updates_1__din),
    .num_updates_out_q_fifo_V_full_n(num_updates_1__full_n),
    .num_updates_out_q_fifo_V_write(num_updates_1__write),
    .update_config_q_fifo_V_dout(update_config_1__dout),
    .update_config_q_fifo_V_empty_n(update_config_1__empty_n),
    .update_config_q_fifo_V_read(update_config_1__read),
    .update_config_q_peek_val(update_config_1__dout),
    .update_out_q_fifo_V_din(update_mm2pe_1__din),
    .update_out_q_fifo_V_full_n(update_mm2pe_1__full_n),
    .update_out_q_fifo_V_write(update_mm2pe_1__write),
    .update_in_q_fifo_V_dout(update_pe2mm_1__dout),
    .update_in_q_fifo_V_empty_n(update_pe2mm_1__empty_n),
    .update_in_q_fifo_V_read(update_pe2mm_1__read),
    .update_in_q_peek_val(update_pe2mm_1__dout),
    .update_phase_q_fifo_V_dout(update_phase_1__dout),
    .update_phase_q_fifo_V_empty_n(update_phase_1__empty_n),
    .update_phase_q_fifo_V_read(update_phase_1__read),
    .update_phase_q_peek_val(update_phase_1__dout),
    .updates_read_addr_q_fifo_V_din(update_read_addr_1__din),
    .updates_read_addr_q_fifo_V_full_n(update_read_addr_1__full_n),
    .updates_read_addr_q_fifo_V_write(update_read_addr_1__write),
    .updates_read_data_q_fifo_V_dout(update_read_data_1__dout),
    .updates_read_data_q_fifo_V_empty_n(update_read_data_1__empty_n),
    .updates_read_data_q_fifo_V_read(update_read_data_1__read),
    .updates_read_data_q_peek_val(update_read_data_1__dout),
    .update_req_q_fifo_V_dout(update_req_1__dout),
    .update_req_q_fifo_V_empty_n(update_req_1__empty_n),
    .update_req_q_fifo_V_read(update_req_1__read),
    .update_req_q_peek_val(update_req_1__dout),
    .updates_write_addr_q_fifo_V_din(update_write_addr_1__din),
    .updates_write_addr_q_fifo_V_full_n(update_write_addr_1__full_n),
    .updates_write_addr_q_fifo_V_write(update_write_addr_1__write),
    .updates_write_data_q_fifo_V_din(update_write_data_1__din),
    .updates_write_data_q_fifo_V_full_n(update_write_data_1__full_n),
    .updates_write_data_q_fifo_V_write(update_write_data_1__write)
  );


  UpdateHandler_UpdateHandler
  UpdateHandler_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateHandler_2__ap_rst_n__q2),
    .ap_start(UpdateHandler_2__ap_start),
    .ap_done(UpdateHandler_2__ap_done),
    .ap_idle(UpdateHandler_2__ap_idle),
    .ap_ready(UpdateHandler_2__ap_ready),
    .num_partitions(UpdateHandler_2___num_partitions__q2),
    .num_updates_out_q_fifo_V_din(num_updates_2__din),
    .num_updates_out_q_fifo_V_full_n(num_updates_2__full_n),
    .num_updates_out_q_fifo_V_write(num_updates_2__write),
    .update_config_q_fifo_V_dout(update_config_2__dout),
    .update_config_q_fifo_V_empty_n(update_config_2__empty_n),
    .update_config_q_fifo_V_read(update_config_2__read),
    .update_config_q_peek_val(update_config_2__dout),
    .update_out_q_fifo_V_din(update_mm2pe_2__din),
    .update_out_q_fifo_V_full_n(update_mm2pe_2__full_n),
    .update_out_q_fifo_V_write(update_mm2pe_2__write),
    .update_in_q_fifo_V_dout(update_pe2mm_2__dout),
    .update_in_q_fifo_V_empty_n(update_pe2mm_2__empty_n),
    .update_in_q_fifo_V_read(update_pe2mm_2__read),
    .update_in_q_peek_val(update_pe2mm_2__dout),
    .update_phase_q_fifo_V_dout(update_phase_2__dout),
    .update_phase_q_fifo_V_empty_n(update_phase_2__empty_n),
    .update_phase_q_fifo_V_read(update_phase_2__read),
    .update_phase_q_peek_val(update_phase_2__dout),
    .updates_read_addr_q_fifo_V_din(update_read_addr_2__din),
    .updates_read_addr_q_fifo_V_full_n(update_read_addr_2__full_n),
    .updates_read_addr_q_fifo_V_write(update_read_addr_2__write),
    .updates_read_data_q_fifo_V_dout(update_read_data_2__dout),
    .updates_read_data_q_fifo_V_empty_n(update_read_data_2__empty_n),
    .updates_read_data_q_fifo_V_read(update_read_data_2__read),
    .updates_read_data_q_peek_val(update_read_data_2__dout),
    .update_req_q_fifo_V_dout(update_req_2__dout),
    .update_req_q_fifo_V_empty_n(update_req_2__empty_n),
    .update_req_q_fifo_V_read(update_req_2__read),
    .update_req_q_peek_val(update_req_2__dout),
    .updates_write_addr_q_fifo_V_din(update_write_addr_2__din),
    .updates_write_addr_q_fifo_V_full_n(update_write_addr_2__full_n),
    .updates_write_addr_q_fifo_V_write(update_write_addr_2__write),
    .updates_write_data_q_fifo_V_din(update_write_data_2__din),
    .updates_write_data_q_fifo_V_full_n(update_write_data_2__full_n),
    .updates_write_data_q_fifo_V_write(update_write_data_2__write)
  );


  UpdateHandler_UpdateHandler
  UpdateHandler_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateHandler_3__ap_rst_n__q2),
    .ap_start(UpdateHandler_3__ap_start),
    .ap_done(UpdateHandler_3__ap_done),
    .ap_idle(UpdateHandler_3__ap_idle),
    .ap_ready(UpdateHandler_3__ap_ready),
    .num_partitions(UpdateHandler_3___num_partitions__q2),
    .num_updates_out_q_fifo_V_din(num_updates_3__din),
    .num_updates_out_q_fifo_V_full_n(num_updates_3__full_n),
    .num_updates_out_q_fifo_V_write(num_updates_3__write),
    .update_config_q_fifo_V_dout(update_config_3__dout),
    .update_config_q_fifo_V_empty_n(update_config_3__empty_n),
    .update_config_q_fifo_V_read(update_config_3__read),
    .update_config_q_peek_val(update_config_3__dout),
    .update_out_q_fifo_V_din(update_mm2pe_3__din),
    .update_out_q_fifo_V_full_n(update_mm2pe_3__full_n),
    .update_out_q_fifo_V_write(update_mm2pe_3__write),
    .update_in_q_fifo_V_dout(update_pe2mm_3__dout),
    .update_in_q_fifo_V_empty_n(update_pe2mm_3__empty_n),
    .update_in_q_fifo_V_read(update_pe2mm_3__read),
    .update_in_q_peek_val(update_pe2mm_3__dout),
    .update_phase_q_fifo_V_dout(update_phase_3__dout),
    .update_phase_q_fifo_V_empty_n(update_phase_3__empty_n),
    .update_phase_q_fifo_V_read(update_phase_3__read),
    .update_phase_q_peek_val(update_phase_3__dout),
    .updates_read_addr_q_fifo_V_din(update_read_addr_3__din),
    .updates_read_addr_q_fifo_V_full_n(update_read_addr_3__full_n),
    .updates_read_addr_q_fifo_V_write(update_read_addr_3__write),
    .updates_read_data_q_fifo_V_dout(update_read_data_3__dout),
    .updates_read_data_q_fifo_V_empty_n(update_read_data_3__empty_n),
    .updates_read_data_q_fifo_V_read(update_read_data_3__read),
    .updates_read_data_q_peek_val(update_read_data_3__dout),
    .update_req_q_fifo_V_dout(update_req_3__dout),
    .update_req_q_fifo_V_empty_n(update_req_3__empty_n),
    .update_req_q_fifo_V_read(update_req_3__read),
    .update_req_q_peek_val(update_req_3__dout),
    .updates_write_addr_q_fifo_V_din(update_write_addr_3__din),
    .updates_write_addr_q_fifo_V_full_n(update_write_addr_3__full_n),
    .updates_write_addr_q_fifo_V_write(update_write_addr_3__write),
    .updates_write_data_q_fifo_V_din(update_write_data_3__din),
    .updates_write_data_q_fifo_V_full_n(update_write_data_3__full_n),
    .updates_write_data_q_fifo_V_write(update_write_data_3__write)
  );


  UpdateHandler_UpdateHandler
  UpdateHandler_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateHandler_4__ap_rst_n__q2),
    .ap_start(UpdateHandler_4__ap_start),
    .ap_done(UpdateHandler_4__ap_done),
    .ap_idle(UpdateHandler_4__ap_idle),
    .ap_ready(UpdateHandler_4__ap_ready),
    .num_partitions(UpdateHandler_4___num_partitions__q2),
    .num_updates_out_q_fifo_V_din(num_updates_4__din),
    .num_updates_out_q_fifo_V_full_n(num_updates_4__full_n),
    .num_updates_out_q_fifo_V_write(num_updates_4__write),
    .update_config_q_fifo_V_dout(update_config_4__dout),
    .update_config_q_fifo_V_empty_n(update_config_4__empty_n),
    .update_config_q_fifo_V_read(update_config_4__read),
    .update_config_q_peek_val(update_config_4__dout),
    .update_out_q_fifo_V_din(update_mm2pe_4__din),
    .update_out_q_fifo_V_full_n(update_mm2pe_4__full_n),
    .update_out_q_fifo_V_write(update_mm2pe_4__write),
    .update_in_q_fifo_V_dout(update_pe2mm_4__dout),
    .update_in_q_fifo_V_empty_n(update_pe2mm_4__empty_n),
    .update_in_q_fifo_V_read(update_pe2mm_4__read),
    .update_in_q_peek_val(update_pe2mm_4__dout),
    .update_phase_q_fifo_V_dout(update_phase_4__dout),
    .update_phase_q_fifo_V_empty_n(update_phase_4__empty_n),
    .update_phase_q_fifo_V_read(update_phase_4__read),
    .update_phase_q_peek_val(update_phase_4__dout),
    .updates_read_addr_q_fifo_V_din(update_read_addr_4__din),
    .updates_read_addr_q_fifo_V_full_n(update_read_addr_4__full_n),
    .updates_read_addr_q_fifo_V_write(update_read_addr_4__write),
    .updates_read_data_q_fifo_V_dout(update_read_data_4__dout),
    .updates_read_data_q_fifo_V_empty_n(update_read_data_4__empty_n),
    .updates_read_data_q_fifo_V_read(update_read_data_4__read),
    .updates_read_data_q_peek_val(update_read_data_4__dout),
    .update_req_q_fifo_V_dout(update_req_4__dout),
    .update_req_q_fifo_V_empty_n(update_req_4__empty_n),
    .update_req_q_fifo_V_read(update_req_4__read),
    .update_req_q_peek_val(update_req_4__dout),
    .updates_write_addr_q_fifo_V_din(update_write_addr_4__din),
    .updates_write_addr_q_fifo_V_full_n(update_write_addr_4__full_n),
    .updates_write_addr_q_fifo_V_write(update_write_addr_4__write),
    .updates_write_data_q_fifo_V_din(update_write_data_4__din),
    .updates_write_data_q_fifo_V_full_n(update_write_data_4__full_n),
    .updates_write_data_q_fifo_V_write(update_write_data_4__write)
  );


  UpdateHandler_UpdateHandler
  UpdateHandler_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateHandler_5__ap_rst_n__q2),
    .ap_start(UpdateHandler_5__ap_start),
    .ap_done(UpdateHandler_5__ap_done),
    .ap_idle(UpdateHandler_5__ap_idle),
    .ap_ready(UpdateHandler_5__ap_ready),
    .num_partitions(UpdateHandler_5___num_partitions__q2),
    .num_updates_out_q_fifo_V_din(num_updates_5__din),
    .num_updates_out_q_fifo_V_full_n(num_updates_5__full_n),
    .num_updates_out_q_fifo_V_write(num_updates_5__write),
    .update_config_q_fifo_V_dout(update_config_5__dout),
    .update_config_q_fifo_V_empty_n(update_config_5__empty_n),
    .update_config_q_fifo_V_read(update_config_5__read),
    .update_config_q_peek_val(update_config_5__dout),
    .update_out_q_fifo_V_din(update_mm2pe_5__din),
    .update_out_q_fifo_V_full_n(update_mm2pe_5__full_n),
    .update_out_q_fifo_V_write(update_mm2pe_5__write),
    .update_in_q_fifo_V_dout(update_pe2mm_5__dout),
    .update_in_q_fifo_V_empty_n(update_pe2mm_5__empty_n),
    .update_in_q_fifo_V_read(update_pe2mm_5__read),
    .update_in_q_peek_val(update_pe2mm_5__dout),
    .update_phase_q_fifo_V_dout(update_phase_5__dout),
    .update_phase_q_fifo_V_empty_n(update_phase_5__empty_n),
    .update_phase_q_fifo_V_read(update_phase_5__read),
    .update_phase_q_peek_val(update_phase_5__dout),
    .updates_read_addr_q_fifo_V_din(update_read_addr_5__din),
    .updates_read_addr_q_fifo_V_full_n(update_read_addr_5__full_n),
    .updates_read_addr_q_fifo_V_write(update_read_addr_5__write),
    .updates_read_data_q_fifo_V_dout(update_read_data_5__dout),
    .updates_read_data_q_fifo_V_empty_n(update_read_data_5__empty_n),
    .updates_read_data_q_fifo_V_read(update_read_data_5__read),
    .updates_read_data_q_peek_val(update_read_data_5__dout),
    .update_req_q_fifo_V_dout(update_req_5__dout),
    .update_req_q_fifo_V_empty_n(update_req_5__empty_n),
    .update_req_q_fifo_V_read(update_req_5__read),
    .update_req_q_peek_val(update_req_5__dout),
    .updates_write_addr_q_fifo_V_din(update_write_addr_5__din),
    .updates_write_addr_q_fifo_V_full_n(update_write_addr_5__full_n),
    .updates_write_addr_q_fifo_V_write(update_write_addr_5__write),
    .updates_write_data_q_fifo_V_din(update_write_data_5__din),
    .updates_write_data_q_fifo_V_full_n(update_write_data_5__full_n),
    .updates_write_data_q_fifo_V_write(update_write_data_5__write)
  );


  UpdateHandler_UpdateHandler
  UpdateHandler_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateHandler_6__ap_rst_n__q2),
    .ap_start(UpdateHandler_6__ap_start),
    .ap_done(UpdateHandler_6__ap_done),
    .ap_idle(UpdateHandler_6__ap_idle),
    .ap_ready(UpdateHandler_6__ap_ready),
    .num_partitions(UpdateHandler_6___num_partitions__q2),
    .num_updates_out_q_fifo_V_din(num_updates_6__din),
    .num_updates_out_q_fifo_V_full_n(num_updates_6__full_n),
    .num_updates_out_q_fifo_V_write(num_updates_6__write),
    .update_config_q_fifo_V_dout(update_config_6__dout),
    .update_config_q_fifo_V_empty_n(update_config_6__empty_n),
    .update_config_q_fifo_V_read(update_config_6__read),
    .update_config_q_peek_val(update_config_6__dout),
    .update_out_q_fifo_V_din(update_mm2pe_6__din),
    .update_out_q_fifo_V_full_n(update_mm2pe_6__full_n),
    .update_out_q_fifo_V_write(update_mm2pe_6__write),
    .update_in_q_fifo_V_dout(update_pe2mm_6__dout),
    .update_in_q_fifo_V_empty_n(update_pe2mm_6__empty_n),
    .update_in_q_fifo_V_read(update_pe2mm_6__read),
    .update_in_q_peek_val(update_pe2mm_6__dout),
    .update_phase_q_fifo_V_dout(update_phase_6__dout),
    .update_phase_q_fifo_V_empty_n(update_phase_6__empty_n),
    .update_phase_q_fifo_V_read(update_phase_6__read),
    .update_phase_q_peek_val(update_phase_6__dout),
    .updates_read_addr_q_fifo_V_din(update_read_addr_6__din),
    .updates_read_addr_q_fifo_V_full_n(update_read_addr_6__full_n),
    .updates_read_addr_q_fifo_V_write(update_read_addr_6__write),
    .updates_read_data_q_fifo_V_dout(update_read_data_6__dout),
    .updates_read_data_q_fifo_V_empty_n(update_read_data_6__empty_n),
    .updates_read_data_q_fifo_V_read(update_read_data_6__read),
    .updates_read_data_q_peek_val(update_read_data_6__dout),
    .update_req_q_fifo_V_dout(update_req_6__dout),
    .update_req_q_fifo_V_empty_n(update_req_6__empty_n),
    .update_req_q_fifo_V_read(update_req_6__read),
    .update_req_q_peek_val(update_req_6__dout),
    .updates_write_addr_q_fifo_V_din(update_write_addr_6__din),
    .updates_write_addr_q_fifo_V_full_n(update_write_addr_6__full_n),
    .updates_write_addr_q_fifo_V_write(update_write_addr_6__write),
    .updates_write_data_q_fifo_V_din(update_write_data_6__din),
    .updates_write_data_q_fifo_V_full_n(update_write_data_6__full_n),
    .updates_write_data_q_fifo_V_write(update_write_data_6__write)
  );


  UpdateHandler_UpdateHandler
  UpdateHandler_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateHandler_7__ap_rst_n__q2),
    .ap_start(UpdateHandler_7__ap_start),
    .ap_done(UpdateHandler_7__ap_done),
    .ap_idle(UpdateHandler_7__ap_idle),
    .ap_ready(UpdateHandler_7__ap_ready),
    .num_partitions(UpdateHandler_7___num_partitions__q2),
    .num_updates_out_q_fifo_V_din(num_updates_7__din),
    .num_updates_out_q_fifo_V_full_n(num_updates_7__full_n),
    .num_updates_out_q_fifo_V_write(num_updates_7__write),
    .update_config_q_fifo_V_dout(update_config_7__dout),
    .update_config_q_fifo_V_empty_n(update_config_7__empty_n),
    .update_config_q_fifo_V_read(update_config_7__read),
    .update_config_q_peek_val(update_config_7__dout),
    .update_out_q_fifo_V_din(update_mm2pe_7__din),
    .update_out_q_fifo_V_full_n(update_mm2pe_7__full_n),
    .update_out_q_fifo_V_write(update_mm2pe_7__write),
    .update_in_q_fifo_V_dout(update_pe2mm_7__dout),
    .update_in_q_fifo_V_empty_n(update_pe2mm_7__empty_n),
    .update_in_q_fifo_V_read(update_pe2mm_7__read),
    .update_in_q_peek_val(update_pe2mm_7__dout),
    .update_phase_q_fifo_V_dout(update_phase_7__dout),
    .update_phase_q_fifo_V_empty_n(update_phase_7__empty_n),
    .update_phase_q_fifo_V_read(update_phase_7__read),
    .update_phase_q_peek_val(update_phase_7__dout),
    .updates_read_addr_q_fifo_V_din(update_read_addr_7__din),
    .updates_read_addr_q_fifo_V_full_n(update_read_addr_7__full_n),
    .updates_read_addr_q_fifo_V_write(update_read_addr_7__write),
    .updates_read_data_q_fifo_V_dout(update_read_data_7__dout),
    .updates_read_data_q_fifo_V_empty_n(update_read_data_7__empty_n),
    .updates_read_data_q_fifo_V_read(update_read_data_7__read),
    .updates_read_data_q_peek_val(update_read_data_7__dout),
    .update_req_q_fifo_V_dout(update_req_7__dout),
    .update_req_q_fifo_V_empty_n(update_req_7__empty_n),
    .update_req_q_fifo_V_read(update_req_7__read),
    .update_req_q_peek_val(update_req_7__dout),
    .updates_write_addr_q_fifo_V_din(update_write_addr_7__din),
    .updates_write_addr_q_fifo_V_full_n(update_write_addr_7__full_n),
    .updates_write_addr_q_fifo_V_write(update_write_addr_7__write),
    .updates_write_data_q_fifo_V_din(update_write_data_7__din),
    .updates_write_data_q_fifo_V_full_n(update_write_data_7__full_n),
    .updates_write_data_q_fifo_V_write(update_write_data_7__write)
  );


  UpdateMem_UpdateMem
  UpdateMem_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateMem_0__ap_rst_n__q2),
    .ap_start(UpdateMem_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .read_addr_q_fifo_V_dout(update_read_addr_0__dout),
    .read_addr_q_fifo_V_empty_n(update_read_addr_0__empty_n),
    .read_addr_q_fifo_V_read(update_read_addr_0__read),
    .read_addr_q_peek_val(update_read_addr_0__dout),
    .read_data_q_fifo_V_din(update_read_data_0__din),
    .read_data_q_fifo_V_full_n(update_read_data_0__full_n),
    .read_data_q_fifo_V_write(update_read_data_0__write),
    .write_addr_q_fifo_V_dout(update_write_addr_0__dout),
    .write_addr_q_fifo_V_empty_n(update_write_addr_0__empty_n),
    .write_addr_q_fifo_V_read(update_write_addr_0__read),
    .write_addr_q_peek_val(update_write_addr_0__dout),
    .write_data_q_fifo_V_dout(update_write_data_0__dout),
    .write_data_q_fifo_V_empty_n(update_write_data_0__empty_n),
    .write_data_q_fifo_V_read(update_write_data_0__read),
    .write_data_q_peek_val(update_write_data_0__dout),
    .updates_read_addr_V_din(updates_0_read_addr__din),
    .updates_read_addr_V_full_n(updates_0_read_addr__full_n),
    .updates_read_addr_V_write(updates_0_read_addr__write),
    .updates_read_data_V_data_V_dout(updates_0_read_data__dout),
    .updates_read_data_V_data_V_empty_n(updates_0_read_data__empty_n),
    .updates_read_data_V_data_V_read(updates_0_read_data__read),
    .updates_write_addr_V_din(updates_0_write_addr__din),
    .updates_write_addr_V_full_n(updates_0_write_addr__full_n),
    .updates_write_addr_V_write(updates_0_write_addr__write),
    .updates_write_data_V_data_V_din(updates_0_write_data__din),
    .updates_write_data_V_data_V_full_n(updates_0_write_data__full_n),
    .updates_write_data_V_data_V_write(updates_0_write_data__write)
  );


  UpdateMem_UpdateMem
  UpdateMem_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateMem_1__ap_rst_n__q2),
    .ap_start(UpdateMem_1__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .read_addr_q_fifo_V_dout(update_read_addr_1__dout),
    .read_addr_q_fifo_V_empty_n(update_read_addr_1__empty_n),
    .read_addr_q_fifo_V_read(update_read_addr_1__read),
    .read_addr_q_peek_val(update_read_addr_1__dout),
    .read_data_q_fifo_V_din(update_read_data_1__din),
    .read_data_q_fifo_V_full_n(update_read_data_1__full_n),
    .read_data_q_fifo_V_write(update_read_data_1__write),
    .write_addr_q_fifo_V_dout(update_write_addr_1__dout),
    .write_addr_q_fifo_V_empty_n(update_write_addr_1__empty_n),
    .write_addr_q_fifo_V_read(update_write_addr_1__read),
    .write_addr_q_peek_val(update_write_addr_1__dout),
    .write_data_q_fifo_V_dout(update_write_data_1__dout),
    .write_data_q_fifo_V_empty_n(update_write_data_1__empty_n),
    .write_data_q_fifo_V_read(update_write_data_1__read),
    .write_data_q_peek_val(update_write_data_1__dout),
    .updates_read_addr_V_din(updates_1_read_addr__din),
    .updates_read_addr_V_full_n(updates_1_read_addr__full_n),
    .updates_read_addr_V_write(updates_1_read_addr__write),
    .updates_read_data_V_data_V_dout(updates_1_read_data__dout),
    .updates_read_data_V_data_V_empty_n(updates_1_read_data__empty_n),
    .updates_read_data_V_data_V_read(updates_1_read_data__read),
    .updates_write_addr_V_din(updates_1_write_addr__din),
    .updates_write_addr_V_full_n(updates_1_write_addr__full_n),
    .updates_write_addr_V_write(updates_1_write_addr__write),
    .updates_write_data_V_data_V_din(updates_1_write_data__din),
    .updates_write_data_V_data_V_full_n(updates_1_write_data__full_n),
    .updates_write_data_V_data_V_write(updates_1_write_data__write)
  );


  UpdateMem_UpdateMem
  UpdateMem_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateMem_2__ap_rst_n__q2),
    .ap_start(UpdateMem_2__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .read_addr_q_fifo_V_dout(update_read_addr_2__dout),
    .read_addr_q_fifo_V_empty_n(update_read_addr_2__empty_n),
    .read_addr_q_fifo_V_read(update_read_addr_2__read),
    .read_addr_q_peek_val(update_read_addr_2__dout),
    .read_data_q_fifo_V_din(update_read_data_2__din),
    .read_data_q_fifo_V_full_n(update_read_data_2__full_n),
    .read_data_q_fifo_V_write(update_read_data_2__write),
    .write_addr_q_fifo_V_dout(update_write_addr_2__dout),
    .write_addr_q_fifo_V_empty_n(update_write_addr_2__empty_n),
    .write_addr_q_fifo_V_read(update_write_addr_2__read),
    .write_addr_q_peek_val(update_write_addr_2__dout),
    .write_data_q_fifo_V_dout(update_write_data_2__dout),
    .write_data_q_fifo_V_empty_n(update_write_data_2__empty_n),
    .write_data_q_fifo_V_read(update_write_data_2__read),
    .write_data_q_peek_val(update_write_data_2__dout),
    .updates_read_addr_V_din(updates_2_read_addr__din),
    .updates_read_addr_V_full_n(updates_2_read_addr__full_n),
    .updates_read_addr_V_write(updates_2_read_addr__write),
    .updates_read_data_V_data_V_dout(updates_2_read_data__dout),
    .updates_read_data_V_data_V_empty_n(updates_2_read_data__empty_n),
    .updates_read_data_V_data_V_read(updates_2_read_data__read),
    .updates_write_addr_V_din(updates_2_write_addr__din),
    .updates_write_addr_V_full_n(updates_2_write_addr__full_n),
    .updates_write_addr_V_write(updates_2_write_addr__write),
    .updates_write_data_V_data_V_din(updates_2_write_data__din),
    .updates_write_data_V_data_V_full_n(updates_2_write_data__full_n),
    .updates_write_data_V_data_V_write(updates_2_write_data__write)
  );


  UpdateMem_UpdateMem
  UpdateMem_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateMem_3__ap_rst_n__q2),
    .ap_start(UpdateMem_3__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .read_addr_q_fifo_V_dout(update_read_addr_3__dout),
    .read_addr_q_fifo_V_empty_n(update_read_addr_3__empty_n),
    .read_addr_q_fifo_V_read(update_read_addr_3__read),
    .read_addr_q_peek_val(update_read_addr_3__dout),
    .read_data_q_fifo_V_din(update_read_data_3__din),
    .read_data_q_fifo_V_full_n(update_read_data_3__full_n),
    .read_data_q_fifo_V_write(update_read_data_3__write),
    .write_addr_q_fifo_V_dout(update_write_addr_3__dout),
    .write_addr_q_fifo_V_empty_n(update_write_addr_3__empty_n),
    .write_addr_q_fifo_V_read(update_write_addr_3__read),
    .write_addr_q_peek_val(update_write_addr_3__dout),
    .write_data_q_fifo_V_dout(update_write_data_3__dout),
    .write_data_q_fifo_V_empty_n(update_write_data_3__empty_n),
    .write_data_q_fifo_V_read(update_write_data_3__read),
    .write_data_q_peek_val(update_write_data_3__dout),
    .updates_read_addr_V_din(updates_3_read_addr__din),
    .updates_read_addr_V_full_n(updates_3_read_addr__full_n),
    .updates_read_addr_V_write(updates_3_read_addr__write),
    .updates_read_data_V_data_V_dout(updates_3_read_data__dout),
    .updates_read_data_V_data_V_empty_n(updates_3_read_data__empty_n),
    .updates_read_data_V_data_V_read(updates_3_read_data__read),
    .updates_write_addr_V_din(updates_3_write_addr__din),
    .updates_write_addr_V_full_n(updates_3_write_addr__full_n),
    .updates_write_addr_V_write(updates_3_write_addr__write),
    .updates_write_data_V_data_V_din(updates_3_write_data__din),
    .updates_write_data_V_data_V_full_n(updates_3_write_data__full_n),
    .updates_write_data_V_data_V_write(updates_3_write_data__write)
  );


  UpdateMem_UpdateMem
  UpdateMem_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateMem_4__ap_rst_n__q2),
    .ap_start(UpdateMem_4__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .read_addr_q_fifo_V_dout(update_read_addr_4__dout),
    .read_addr_q_fifo_V_empty_n(update_read_addr_4__empty_n),
    .read_addr_q_fifo_V_read(update_read_addr_4__read),
    .read_addr_q_peek_val(update_read_addr_4__dout),
    .read_data_q_fifo_V_din(update_read_data_4__din),
    .read_data_q_fifo_V_full_n(update_read_data_4__full_n),
    .read_data_q_fifo_V_write(update_read_data_4__write),
    .write_addr_q_fifo_V_dout(update_write_addr_4__dout),
    .write_addr_q_fifo_V_empty_n(update_write_addr_4__empty_n),
    .write_addr_q_fifo_V_read(update_write_addr_4__read),
    .write_addr_q_peek_val(update_write_addr_4__dout),
    .write_data_q_fifo_V_dout(update_write_data_4__dout),
    .write_data_q_fifo_V_empty_n(update_write_data_4__empty_n),
    .write_data_q_fifo_V_read(update_write_data_4__read),
    .write_data_q_peek_val(update_write_data_4__dout),
    .updates_read_addr_V_din(updates_4_read_addr__din),
    .updates_read_addr_V_full_n(updates_4_read_addr__full_n),
    .updates_read_addr_V_write(updates_4_read_addr__write),
    .updates_read_data_V_data_V_dout(updates_4_read_data__dout),
    .updates_read_data_V_data_V_empty_n(updates_4_read_data__empty_n),
    .updates_read_data_V_data_V_read(updates_4_read_data__read),
    .updates_write_addr_V_din(updates_4_write_addr__din),
    .updates_write_addr_V_full_n(updates_4_write_addr__full_n),
    .updates_write_addr_V_write(updates_4_write_addr__write),
    .updates_write_data_V_data_V_din(updates_4_write_data__din),
    .updates_write_data_V_data_V_full_n(updates_4_write_data__full_n),
    .updates_write_data_V_data_V_write(updates_4_write_data__write)
  );


  UpdateMem_UpdateMem
  UpdateMem_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateMem_5__ap_rst_n__q2),
    .ap_start(UpdateMem_5__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .read_addr_q_fifo_V_dout(update_read_addr_5__dout),
    .read_addr_q_fifo_V_empty_n(update_read_addr_5__empty_n),
    .read_addr_q_fifo_V_read(update_read_addr_5__read),
    .read_addr_q_peek_val(update_read_addr_5__dout),
    .read_data_q_fifo_V_din(update_read_data_5__din),
    .read_data_q_fifo_V_full_n(update_read_data_5__full_n),
    .read_data_q_fifo_V_write(update_read_data_5__write),
    .write_addr_q_fifo_V_dout(update_write_addr_5__dout),
    .write_addr_q_fifo_V_empty_n(update_write_addr_5__empty_n),
    .write_addr_q_fifo_V_read(update_write_addr_5__read),
    .write_addr_q_peek_val(update_write_addr_5__dout),
    .write_data_q_fifo_V_dout(update_write_data_5__dout),
    .write_data_q_fifo_V_empty_n(update_write_data_5__empty_n),
    .write_data_q_fifo_V_read(update_write_data_5__read),
    .write_data_q_peek_val(update_write_data_5__dout),
    .updates_read_addr_V_din(updates_5_read_addr__din),
    .updates_read_addr_V_full_n(updates_5_read_addr__full_n),
    .updates_read_addr_V_write(updates_5_read_addr__write),
    .updates_read_data_V_data_V_dout(updates_5_read_data__dout),
    .updates_read_data_V_data_V_empty_n(updates_5_read_data__empty_n),
    .updates_read_data_V_data_V_read(updates_5_read_data__read),
    .updates_write_addr_V_din(updates_5_write_addr__din),
    .updates_write_addr_V_full_n(updates_5_write_addr__full_n),
    .updates_write_addr_V_write(updates_5_write_addr__write),
    .updates_write_data_V_data_V_din(updates_5_write_data__din),
    .updates_write_data_V_data_V_full_n(updates_5_write_data__full_n),
    .updates_write_data_V_data_V_write(updates_5_write_data__write)
  );


  UpdateMem_UpdateMem
  UpdateMem_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateMem_6__ap_rst_n__q2),
    .ap_start(UpdateMem_6__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .read_addr_q_fifo_V_dout(update_read_addr_6__dout),
    .read_addr_q_fifo_V_empty_n(update_read_addr_6__empty_n),
    .read_addr_q_fifo_V_read(update_read_addr_6__read),
    .read_addr_q_peek_val(update_read_addr_6__dout),
    .read_data_q_fifo_V_din(update_read_data_6__din),
    .read_data_q_fifo_V_full_n(update_read_data_6__full_n),
    .read_data_q_fifo_V_write(update_read_data_6__write),
    .write_addr_q_fifo_V_dout(update_write_addr_6__dout),
    .write_addr_q_fifo_V_empty_n(update_write_addr_6__empty_n),
    .write_addr_q_fifo_V_read(update_write_addr_6__read),
    .write_addr_q_peek_val(update_write_addr_6__dout),
    .write_data_q_fifo_V_dout(update_write_data_6__dout),
    .write_data_q_fifo_V_empty_n(update_write_data_6__empty_n),
    .write_data_q_fifo_V_read(update_write_data_6__read),
    .write_data_q_peek_val(update_write_data_6__dout),
    .updates_read_addr_V_din(updates_6_read_addr__din),
    .updates_read_addr_V_full_n(updates_6_read_addr__full_n),
    .updates_read_addr_V_write(updates_6_read_addr__write),
    .updates_read_data_V_data_V_dout(updates_6_read_data__dout),
    .updates_read_data_V_data_V_empty_n(updates_6_read_data__empty_n),
    .updates_read_data_V_data_V_read(updates_6_read_data__read),
    .updates_write_addr_V_din(updates_6_write_addr__din),
    .updates_write_addr_V_full_n(updates_6_write_addr__full_n),
    .updates_write_addr_V_write(updates_6_write_addr__write),
    .updates_write_data_V_data_V_din(updates_6_write_data__din),
    .updates_write_data_V_data_V_full_n(updates_6_write_data__full_n),
    .updates_write_data_V_data_V_write(updates_6_write_data__write)
  );


  UpdateMem_UpdateMem
  UpdateMem_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(UpdateMem_7__ap_rst_n__q2),
    .ap_start(UpdateMem_7__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .read_addr_q_fifo_V_dout(update_read_addr_7__dout),
    .read_addr_q_fifo_V_empty_n(update_read_addr_7__empty_n),
    .read_addr_q_fifo_V_read(update_read_addr_7__read),
    .read_addr_q_peek_val(update_read_addr_7__dout),
    .read_data_q_fifo_V_din(update_read_data_7__din),
    .read_data_q_fifo_V_full_n(update_read_data_7__full_n),
    .read_data_q_fifo_V_write(update_read_data_7__write),
    .write_addr_q_fifo_V_dout(update_write_addr_7__dout),
    .write_addr_q_fifo_V_empty_n(update_write_addr_7__empty_n),
    .write_addr_q_fifo_V_read(update_write_addr_7__read),
    .write_addr_q_peek_val(update_write_addr_7__dout),
    .write_data_q_fifo_V_dout(update_write_data_7__dout),
    .write_data_q_fifo_V_empty_n(update_write_data_7__empty_n),
    .write_data_q_fifo_V_read(update_write_data_7__read),
    .write_data_q_peek_val(update_write_data_7__dout),
    .updates_read_addr_V_din(updates_7_read_addr__din),
    .updates_read_addr_V_full_n(updates_7_read_addr__full_n),
    .updates_read_addr_V_write(updates_7_read_addr__write),
    .updates_read_data_V_data_V_dout(updates_7_read_data__dout),
    .updates_read_data_V_data_V_empty_n(updates_7_read_data__empty_n),
    .updates_read_data_V_data_V_read(updates_7_read_data__read),
    .updates_write_addr_V_din(updates_7_write_addr__din),
    .updates_write_addr_V_full_n(updates_7_write_addr__full_n),
    .updates_write_addr_V_write(updates_7_write_addr__write),
    .updates_write_data_V_data_V_din(updates_7_write_data__din),
    .updates_write_data_V_data_V_full_n(updates_7_write_data__full_n),
    .updates_write_data_V_data_V_write(updates_7_write_data__write)
  );


  VertexMem_VertexMem
  VertexMem_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(VertexMem_0__ap_rst_n__q2),
    .ap_start(VertexMem_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .degrees_read_addr_V_din(degrees_read_addr__din),
    .degrees_read_addr_V_full_n(degrees_read_addr__full_n),
    .degrees_read_addr_V_write(degrees_read_addr__write),
    .degrees_read_data_V_data_V_dout(degrees_read_data__dout),
    .degrees_read_data_V_data_V_empty_n(degrees_read_data__empty_n),
    .degrees_read_data_V_data_V_read(degrees_read_data__read),
    .rankings_read_addr_V_din(rankings_read_addr__din),
    .rankings_read_addr_V_full_n(rankings_read_addr__full_n),
    .rankings_read_addr_V_write(rankings_read_addr__write),
    .rankings_read_data_V_data_V_dout(rankings_read_data__dout),
    .rankings_read_data_V_data_V_empty_n(rankings_read_data__empty_n),
    .rankings_read_data_V_data_V_read(rankings_read_data__read),
    .rankings_write_addr_V_din(rankings_write_addr__din),
    .rankings_write_addr_V_full_n(rankings_write_addr__full_n),
    .rankings_write_addr_V_write(rankings_write_addr__write),
    .rankings_write_data_V_data_V_din(rankings_write_data__din),
    .rankings_write_data_V_data_V_full_n(rankings_write_data__full_n),
    .rankings_write_data_V_data_V_write(rankings_write_data__write),
    .scatter_req_q_fifo_V_dout(scatter_phase_vertex_req__dout),
    .scatter_req_q_fifo_V_empty_n(scatter_phase_vertex_req__empty_n),
    .scatter_req_q_fifo_V_read(scatter_phase_vertex_req__read),
    .scatter_req_q_peek_val(scatter_phase_vertex_req__dout),
    .tmps_read_addr_V_din(tmps_read_addr__din),
    .tmps_read_addr_V_full_n(tmps_read_addr__full_n),
    .tmps_read_addr_V_write(tmps_read_addr__write),
    .tmps_read_data_V_data_V_dout(tmps_read_data__dout),
    .tmps_read_data_V_data_V_empty_n(tmps_read_data__empty_n),
    .tmps_read_data_V_data_V_read(tmps_read_data__read),
    .tmps_write_addr_V_din(tmps_write_addr__din),
    .tmps_write_addr_V_full_n(tmps_write_addr__full_n),
    .tmps_write_addr_V_write(tmps_write_addr__write),
    .tmps_write_data_V_data_V_din(tmps_write_data__din),
    .tmps_write_data_V_data_V_full_n(tmps_write_data__full_n),
    .tmps_write_data_V_data_V_write(tmps_write_data__write),
    .vertex_out_q_fifo_V_0_din(vertex_mm2pe_r0_0__din),
    .vertex_out_q_fifo_V_0_full_n(vertex_mm2pe_r0_0__full_n),
    .vertex_out_q_fifo_V_0_write(vertex_mm2pe_r0_0__write),
    .vertex_out_q_fifo_V_1_din(vertex_mm2pe_r0_1__din),
    .vertex_out_q_fifo_V_1_full_n(vertex_mm2pe_r0_1__full_n),
    .vertex_out_q_fifo_V_1_write(vertex_mm2pe_r0_1__write),
    .vertex_in_q_fifo_V_0_dout(vertex_pe2mm_r0_0__dout),
    .vertex_in_q_fifo_V_0_empty_n(vertex_pe2mm_r0_0__empty_n),
    .vertex_in_q_fifo_V_0_read(vertex_pe2mm_r0_0__read),
    .vertex_in_q_peek_val_0(vertex_pe2mm_r0_0__dout),
    .vertex_in_q_fifo_V_1_dout(vertex_pe2mm_r0_1__dout),
    .vertex_in_q_fifo_V_1_empty_n(vertex_pe2mm_r0_1__empty_n),
    .vertex_in_q_fifo_V_1_read(vertex_pe2mm_r0_1__read),
    .vertex_in_q_peek_val_1(vertex_pe2mm_r0_1__dout),
    .vertex_req_q_fifo_V_0_dout(vertex_req_r0_0__dout),
    .vertex_req_q_fifo_V_0_empty_n(vertex_req_r0_0__empty_n),
    .vertex_req_q_fifo_V_0_read(vertex_req_r0_0__read),
    .vertex_req_q_peek_val_0(vertex_req_r0_0__dout),
    .vertex_req_q_fifo_V_1_dout(vertex_req_r0_1__dout),
    .vertex_req_q_fifo_V_1_empty_n(vertex_req_r0_1__empty_n),
    .vertex_req_q_fifo_V_1_read(vertex_req_r0_1__read),
    .vertex_req_q_peek_val_1(vertex_req_r0_1__dout)
  );


  VertexRouterR1_VertexRouterR1
  VertexRouterR1_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(VertexRouterR1_0__ap_rst_n__q2),
    .ap_start(VertexRouterR1_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .mm_in_q_fifo_V_dout(vertex_mm2pe_r0_1__dout),
    .mm_in_q_fifo_V_empty_n(vertex_mm2pe_r0_1__empty_n),
    .mm_in_q_fifo_V_read(vertex_mm2pe_r0_1__read),
    .pe_out_q_fifo_V_0_din(vertex_mm2pe_r1_0__din),
    .pe_out_q_fifo_V_0_full_n(vertex_mm2pe_r1_0__full_n),
    .pe_out_q_fifo_V_0_write(vertex_mm2pe_r1_0__write),
    .pe_out_q_fifo_V_1_din(vertex_mm2pe_r1_1__din),
    .pe_out_q_fifo_V_1_full_n(vertex_mm2pe_r1_1__full_n),
    .pe_out_q_fifo_V_1_write(vertex_mm2pe_r1_1__write),
    .pe_out_q_fifo_V_2_din(vertex_mm2pe_r1_2__din),
    .pe_out_q_fifo_V_2_full_n(vertex_mm2pe_r1_2__full_n),
    .pe_out_q_fifo_V_2_write(vertex_mm2pe_r1_2__write),
    .pe_out_q_fifo_V_3_din(vertex_mm2pe_r1_3__din),
    .pe_out_q_fifo_V_3_full_n(vertex_mm2pe_r1_3__full_n),
    .pe_out_q_fifo_V_3_write(vertex_mm2pe_r1_3__write),
    .mm_out_q_fifo_V_din(vertex_pe2mm_r0_1__din),
    .mm_out_q_fifo_V_full_n(vertex_pe2mm_r0_1__full_n),
    .mm_out_q_fifo_V_write(vertex_pe2mm_r0_1__write),
    .pe_in_q_fifo_V_0_dout(vertex_pe2mm_r1_0__dout),
    .pe_in_q_fifo_V_0_empty_n(vertex_pe2mm_r1_0__empty_n),
    .pe_in_q_fifo_V_0_read(vertex_pe2mm_r1_0__read),
    .pe_in_q_peek_val_0(vertex_pe2mm_r1_0__dout),
    .pe_in_q_fifo_V_1_dout(vertex_pe2mm_r1_1__dout),
    .pe_in_q_fifo_V_1_empty_n(vertex_pe2mm_r1_1__empty_n),
    .pe_in_q_fifo_V_1_read(vertex_pe2mm_r1_1__read),
    .pe_in_q_peek_val_1(vertex_pe2mm_r1_1__dout),
    .pe_in_q_fifo_V_2_dout(vertex_pe2mm_r1_2__dout),
    .pe_in_q_fifo_V_2_empty_n(vertex_pe2mm_r1_2__empty_n),
    .pe_in_q_fifo_V_2_read(vertex_pe2mm_r1_2__read),
    .pe_in_q_peek_val_2(vertex_pe2mm_r1_2__dout),
    .pe_in_q_fifo_V_3_dout(vertex_pe2mm_r1_3__dout),
    .pe_in_q_fifo_V_3_empty_n(vertex_pe2mm_r1_3__empty_n),
    .pe_in_q_fifo_V_3_read(vertex_pe2mm_r1_3__read),
    .pe_in_q_peek_val_3(vertex_pe2mm_r1_3__dout),
    .mm_req_q_fifo_V_din(vertex_req_r0_1__din),
    .mm_req_q_fifo_V_full_n(vertex_req_r0_1__full_n),
    .mm_req_q_fifo_V_write(vertex_req_r0_1__write),
    .pe_req_q_fifo_V_0_dout(vertex_req_r1_0__dout),
    .pe_req_q_fifo_V_0_empty_n(vertex_req_r1_0__empty_n),
    .pe_req_q_fifo_V_0_read(vertex_req_r1_0__read),
    .pe_req_q_peek_val_0(vertex_req_r1_0__dout),
    .pe_req_q_fifo_V_1_dout(vertex_req_r1_1__dout),
    .pe_req_q_fifo_V_1_empty_n(vertex_req_r1_1__empty_n),
    .pe_req_q_fifo_V_1_read(vertex_req_r1_1__read),
    .pe_req_q_peek_val_1(vertex_req_r1_1__dout),
    .pe_req_q_fifo_V_2_dout(vertex_req_r1_2__dout),
    .pe_req_q_fifo_V_2_empty_n(vertex_req_r1_2__empty_n),
    .pe_req_q_fifo_V_2_read(vertex_req_r1_2__read),
    .pe_req_q_peek_val_2(vertex_req_r1_2__dout),
    .pe_req_q_fifo_V_3_dout(vertex_req_r1_3__dout),
    .pe_req_q_fifo_V_3_empty_n(vertex_req_r1_3__empty_n),
    .pe_req_q_fifo_V_3_read(vertex_req_r1_3__read),
    .pe_req_q_peek_val_3(vertex_req_r1_3__dout)
  );


  VertexRouterR2_VertexRouterR2
  VertexRouterR2_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(VertexRouterR2_0__ap_rst_n__q2),
    .ap_start(VertexRouterR2_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .mm_in_q_fifo_V_dout(vertex_mm2pe_r1_3__dout),
    .mm_in_q_fifo_V_empty_n(vertex_mm2pe_r1_3__empty_n),
    .mm_in_q_fifo_V_read(vertex_mm2pe_r1_3__read),
    .pe_out_q_fifo_V_0_din(vertex_mm2pe_r2_0__din),
    .pe_out_q_fifo_V_0_full_n(vertex_mm2pe_r2_0__full_n),
    .pe_out_q_fifo_V_0_write(vertex_mm2pe_r2_0__write),
    .pe_out_q_fifo_V_1_din(vertex_mm2pe_r2_1__din),
    .pe_out_q_fifo_V_1_full_n(vertex_mm2pe_r2_1__full_n),
    .pe_out_q_fifo_V_1_write(vertex_mm2pe_r2_1__write),
    .pe_out_q_fifo_V_2_din(vertex_mm2pe_r2_2__din),
    .pe_out_q_fifo_V_2_full_n(vertex_mm2pe_r2_2__full_n),
    .pe_out_q_fifo_V_2_write(vertex_mm2pe_r2_2__write),
    .pe_out_q_fifo_V_3_din(vertex_mm2pe_r2_3__din),
    .pe_out_q_fifo_V_3_full_n(vertex_mm2pe_r2_3__full_n),
    .pe_out_q_fifo_V_3_write(vertex_mm2pe_r2_3__write),
    .mm_out_q_fifo_V_din(vertex_pe2mm_r1_3__din),
    .mm_out_q_fifo_V_full_n(vertex_pe2mm_r1_3__full_n),
    .mm_out_q_fifo_V_write(vertex_pe2mm_r1_3__write),
    .pe_in_q_fifo_V_0_dout(vertex_pe2mm_r2_0__dout),
    .pe_in_q_fifo_V_0_empty_n(vertex_pe2mm_r2_0__empty_n),
    .pe_in_q_fifo_V_0_read(vertex_pe2mm_r2_0__read),
    .pe_in_q_peek_val_0(vertex_pe2mm_r2_0__dout),
    .pe_in_q_fifo_V_1_dout(vertex_pe2mm_r2_1__dout),
    .pe_in_q_fifo_V_1_empty_n(vertex_pe2mm_r2_1__empty_n),
    .pe_in_q_fifo_V_1_read(vertex_pe2mm_r2_1__read),
    .pe_in_q_peek_val_1(vertex_pe2mm_r2_1__dout),
    .pe_in_q_fifo_V_2_dout(vertex_pe2mm_r2_2__dout),
    .pe_in_q_fifo_V_2_empty_n(vertex_pe2mm_r2_2__empty_n),
    .pe_in_q_fifo_V_2_read(vertex_pe2mm_r2_2__read),
    .pe_in_q_peek_val_2(vertex_pe2mm_r2_2__dout),
    .pe_in_q_fifo_V_3_dout(vertex_pe2mm_r2_3__dout),
    .pe_in_q_fifo_V_3_empty_n(vertex_pe2mm_r2_3__empty_n),
    .pe_in_q_fifo_V_3_read(vertex_pe2mm_r2_3__read),
    .pe_in_q_peek_val_3(vertex_pe2mm_r2_3__dout),
    .mm_req_q_fifo_V_din(vertex_req_r1_3__din),
    .mm_req_q_fifo_V_full_n(vertex_req_r1_3__full_n),
    .mm_req_q_fifo_V_write(vertex_req_r1_3__write),
    .pe_req_q_fifo_V_0_dout(vertex_req_r2_0__dout),
    .pe_req_q_fifo_V_0_empty_n(vertex_req_r2_0__empty_n),
    .pe_req_q_fifo_V_0_read(vertex_req_r2_0__read),
    .pe_req_q_peek_val_0(vertex_req_r2_0__dout),
    .pe_req_q_fifo_V_1_dout(vertex_req_r2_1__dout),
    .pe_req_q_fifo_V_1_empty_n(vertex_req_r2_1__empty_n),
    .pe_req_q_fifo_V_1_read(vertex_req_r2_1__read),
    .pe_req_q_peek_val_1(vertex_req_r2_1__dout),
    .pe_req_q_fifo_V_2_dout(vertex_req_r2_2__dout),
    .pe_req_q_fifo_V_2_empty_n(vertex_req_r2_2__empty_n),
    .pe_req_q_fifo_V_2_read(vertex_req_r2_2__read),
    .pe_req_q_peek_val_2(vertex_req_r2_2__dout),
    .pe_req_q_fifo_V_3_dout(vertex_req_r2_3__dout),
    .pe_req_q_fifo_V_3_empty_n(vertex_req_r2_3__empty_n),
    .pe_req_q_fifo_V_3_read(vertex_req_r2_3__read),
    .pe_req_q_peek_val_3(vertex_req_r2_3__dout)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  edges_0__m_axi
  (
    .clk(ap_clk),
    .rst(edges_0__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_edges_0_ARADDR),
    .m_axi_ARBURST(m_axi_edges_0_ARBURST),
    .m_axi_ARCACHE(m_axi_edges_0_ARCACHE),
    .m_axi_ARID(m_axi_edges_0_ARID),
    .m_axi_ARLEN(m_axi_edges_0_ARLEN),
    .m_axi_ARLOCK(m_axi_edges_0_ARLOCK),
    .m_axi_ARPROT(m_axi_edges_0_ARPROT),
    .m_axi_ARQOS(m_axi_edges_0_ARQOS),
    .m_axi_ARREADY(m_axi_edges_0_ARREADY),
    .m_axi_ARREGION(m_axi_edges_0_ARREGION),
    .m_axi_ARSIZE(m_axi_edges_0_ARSIZE),
    .m_axi_ARUSER(m_axi_edges_0_ARUSER),
    .m_axi_ARVALID(m_axi_edges_0_ARVALID),
    .m_axi_AWADDR(m_axi_edges_0_AWADDR),
    .m_axi_AWBURST(m_axi_edges_0_AWBURST),
    .m_axi_AWCACHE(m_axi_edges_0_AWCACHE),
    .m_axi_AWID(m_axi_edges_0_AWID),
    .m_axi_AWLEN(m_axi_edges_0_AWLEN),
    .m_axi_AWLOCK(m_axi_edges_0_AWLOCK),
    .m_axi_AWPROT(m_axi_edges_0_AWPROT),
    .m_axi_AWQOS(m_axi_edges_0_AWQOS),
    .m_axi_AWREADY(m_axi_edges_0_AWREADY),
    .m_axi_AWREGION(m_axi_edges_0_AWREGION),
    .m_axi_AWSIZE(m_axi_edges_0_AWSIZE),
    .m_axi_AWUSER(m_axi_edges_0_AWUSER),
    .m_axi_AWVALID(m_axi_edges_0_AWVALID),
    .m_axi_BID(m_axi_edges_0_BID),
    .m_axi_BREADY(m_axi_edges_0_BREADY),
    .m_axi_BRESP(m_axi_edges_0_BRESP),
    .m_axi_BUSER(m_axi_edges_0_BUSER),
    .m_axi_BVALID(m_axi_edges_0_BVALID),
    .m_axi_RDATA(m_axi_edges_0_RDATA),
    .m_axi_RID(m_axi_edges_0_RID),
    .m_axi_RLAST(m_axi_edges_0_RLAST),
    .m_axi_RREADY(m_axi_edges_0_RREADY),
    .m_axi_RRESP(m_axi_edges_0_RRESP),
    .m_axi_RUSER(m_axi_edges_0_RUSER),
    .m_axi_RVALID(m_axi_edges_0_RVALID),
    .m_axi_WDATA(m_axi_edges_0_WDATA),
    .m_axi_WID(m_axi_edges_0_WID),
    .m_axi_WLAST(m_axi_edges_0_WLAST),
    .m_axi_WREADY(m_axi_edges_0_WREADY),
    .m_axi_WSTRB(m_axi_edges_0_WSTRB),
    .m_axi_WUSER(m_axi_edges_0_WUSER),
    .m_axi_WVALID(m_axi_edges_0_WVALID),
    .read_addr_din(edges_0__q2 + {edges_0_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(edges_0_read_addr__full_n),
    .read_addr_write(edges_0_read_addr__write),
    .read_data_dout(edges_0_read_data__dout),
    .read_data_empty_n(edges_0_read_data__empty_n),
    .read_data_read(edges_0_read_data__read),
    .write_addr_din('d0),
    .write_addr_full_n(),
    .write_addr_write(1'b0),
    .write_data_din('d0),
    .write_data_full_n(),
    .write_data_write(1'b0)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  edges_1__m_axi
  (
    .clk(ap_clk),
    .rst(edges_1__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_edges_1_ARADDR),
    .m_axi_ARBURST(m_axi_edges_1_ARBURST),
    .m_axi_ARCACHE(m_axi_edges_1_ARCACHE),
    .m_axi_ARID(m_axi_edges_1_ARID),
    .m_axi_ARLEN(m_axi_edges_1_ARLEN),
    .m_axi_ARLOCK(m_axi_edges_1_ARLOCK),
    .m_axi_ARPROT(m_axi_edges_1_ARPROT),
    .m_axi_ARQOS(m_axi_edges_1_ARQOS),
    .m_axi_ARREADY(m_axi_edges_1_ARREADY),
    .m_axi_ARREGION(m_axi_edges_1_ARREGION),
    .m_axi_ARSIZE(m_axi_edges_1_ARSIZE),
    .m_axi_ARUSER(m_axi_edges_1_ARUSER),
    .m_axi_ARVALID(m_axi_edges_1_ARVALID),
    .m_axi_AWADDR(m_axi_edges_1_AWADDR),
    .m_axi_AWBURST(m_axi_edges_1_AWBURST),
    .m_axi_AWCACHE(m_axi_edges_1_AWCACHE),
    .m_axi_AWID(m_axi_edges_1_AWID),
    .m_axi_AWLEN(m_axi_edges_1_AWLEN),
    .m_axi_AWLOCK(m_axi_edges_1_AWLOCK),
    .m_axi_AWPROT(m_axi_edges_1_AWPROT),
    .m_axi_AWQOS(m_axi_edges_1_AWQOS),
    .m_axi_AWREADY(m_axi_edges_1_AWREADY),
    .m_axi_AWREGION(m_axi_edges_1_AWREGION),
    .m_axi_AWSIZE(m_axi_edges_1_AWSIZE),
    .m_axi_AWUSER(m_axi_edges_1_AWUSER),
    .m_axi_AWVALID(m_axi_edges_1_AWVALID),
    .m_axi_BID(m_axi_edges_1_BID),
    .m_axi_BREADY(m_axi_edges_1_BREADY),
    .m_axi_BRESP(m_axi_edges_1_BRESP),
    .m_axi_BUSER(m_axi_edges_1_BUSER),
    .m_axi_BVALID(m_axi_edges_1_BVALID),
    .m_axi_RDATA(m_axi_edges_1_RDATA),
    .m_axi_RID(m_axi_edges_1_RID),
    .m_axi_RLAST(m_axi_edges_1_RLAST),
    .m_axi_RREADY(m_axi_edges_1_RREADY),
    .m_axi_RRESP(m_axi_edges_1_RRESP),
    .m_axi_RUSER(m_axi_edges_1_RUSER),
    .m_axi_RVALID(m_axi_edges_1_RVALID),
    .m_axi_WDATA(m_axi_edges_1_WDATA),
    .m_axi_WID(m_axi_edges_1_WID),
    .m_axi_WLAST(m_axi_edges_1_WLAST),
    .m_axi_WREADY(m_axi_edges_1_WREADY),
    .m_axi_WSTRB(m_axi_edges_1_WSTRB),
    .m_axi_WUSER(m_axi_edges_1_WUSER),
    .m_axi_WVALID(m_axi_edges_1_WVALID),
    .read_addr_din(edges_1__q2 + {edges_1_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(edges_1_read_addr__full_n),
    .read_addr_write(edges_1_read_addr__write),
    .read_data_dout(edges_1_read_data__dout),
    .read_data_empty_n(edges_1_read_data__empty_n),
    .read_data_read(edges_1_read_data__read),
    .write_addr_din('d0),
    .write_addr_full_n(),
    .write_addr_write(1'b0),
    .write_data_din('d0),
    .write_data_full_n(),
    .write_data_write(1'b0)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  edges_2__m_axi
  (
    .clk(ap_clk),
    .rst(edges_2__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_edges_2_ARADDR),
    .m_axi_ARBURST(m_axi_edges_2_ARBURST),
    .m_axi_ARCACHE(m_axi_edges_2_ARCACHE),
    .m_axi_ARID(m_axi_edges_2_ARID),
    .m_axi_ARLEN(m_axi_edges_2_ARLEN),
    .m_axi_ARLOCK(m_axi_edges_2_ARLOCK),
    .m_axi_ARPROT(m_axi_edges_2_ARPROT),
    .m_axi_ARQOS(m_axi_edges_2_ARQOS),
    .m_axi_ARREADY(m_axi_edges_2_ARREADY),
    .m_axi_ARREGION(m_axi_edges_2_ARREGION),
    .m_axi_ARSIZE(m_axi_edges_2_ARSIZE),
    .m_axi_ARUSER(m_axi_edges_2_ARUSER),
    .m_axi_ARVALID(m_axi_edges_2_ARVALID),
    .m_axi_AWADDR(m_axi_edges_2_AWADDR),
    .m_axi_AWBURST(m_axi_edges_2_AWBURST),
    .m_axi_AWCACHE(m_axi_edges_2_AWCACHE),
    .m_axi_AWID(m_axi_edges_2_AWID),
    .m_axi_AWLEN(m_axi_edges_2_AWLEN),
    .m_axi_AWLOCK(m_axi_edges_2_AWLOCK),
    .m_axi_AWPROT(m_axi_edges_2_AWPROT),
    .m_axi_AWQOS(m_axi_edges_2_AWQOS),
    .m_axi_AWREADY(m_axi_edges_2_AWREADY),
    .m_axi_AWREGION(m_axi_edges_2_AWREGION),
    .m_axi_AWSIZE(m_axi_edges_2_AWSIZE),
    .m_axi_AWUSER(m_axi_edges_2_AWUSER),
    .m_axi_AWVALID(m_axi_edges_2_AWVALID),
    .m_axi_BID(m_axi_edges_2_BID),
    .m_axi_BREADY(m_axi_edges_2_BREADY),
    .m_axi_BRESP(m_axi_edges_2_BRESP),
    .m_axi_BUSER(m_axi_edges_2_BUSER),
    .m_axi_BVALID(m_axi_edges_2_BVALID),
    .m_axi_RDATA(m_axi_edges_2_RDATA),
    .m_axi_RID(m_axi_edges_2_RID),
    .m_axi_RLAST(m_axi_edges_2_RLAST),
    .m_axi_RREADY(m_axi_edges_2_RREADY),
    .m_axi_RRESP(m_axi_edges_2_RRESP),
    .m_axi_RUSER(m_axi_edges_2_RUSER),
    .m_axi_RVALID(m_axi_edges_2_RVALID),
    .m_axi_WDATA(m_axi_edges_2_WDATA),
    .m_axi_WID(m_axi_edges_2_WID),
    .m_axi_WLAST(m_axi_edges_2_WLAST),
    .m_axi_WREADY(m_axi_edges_2_WREADY),
    .m_axi_WSTRB(m_axi_edges_2_WSTRB),
    .m_axi_WUSER(m_axi_edges_2_WUSER),
    .m_axi_WVALID(m_axi_edges_2_WVALID),
    .read_addr_din(edges_2__q2 + {edges_2_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(edges_2_read_addr__full_n),
    .read_addr_write(edges_2_read_addr__write),
    .read_data_dout(edges_2_read_data__dout),
    .read_data_empty_n(edges_2_read_data__empty_n),
    .read_data_read(edges_2_read_data__read),
    .write_addr_din('d0),
    .write_addr_full_n(),
    .write_addr_write(1'b0),
    .write_data_din('d0),
    .write_data_full_n(),
    .write_data_write(1'b0)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  edges_3__m_axi
  (
    .clk(ap_clk),
    .rst(edges_3__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_edges_3_ARADDR),
    .m_axi_ARBURST(m_axi_edges_3_ARBURST),
    .m_axi_ARCACHE(m_axi_edges_3_ARCACHE),
    .m_axi_ARID(m_axi_edges_3_ARID),
    .m_axi_ARLEN(m_axi_edges_3_ARLEN),
    .m_axi_ARLOCK(m_axi_edges_3_ARLOCK),
    .m_axi_ARPROT(m_axi_edges_3_ARPROT),
    .m_axi_ARQOS(m_axi_edges_3_ARQOS),
    .m_axi_ARREADY(m_axi_edges_3_ARREADY),
    .m_axi_ARREGION(m_axi_edges_3_ARREGION),
    .m_axi_ARSIZE(m_axi_edges_3_ARSIZE),
    .m_axi_ARUSER(m_axi_edges_3_ARUSER),
    .m_axi_ARVALID(m_axi_edges_3_ARVALID),
    .m_axi_AWADDR(m_axi_edges_3_AWADDR),
    .m_axi_AWBURST(m_axi_edges_3_AWBURST),
    .m_axi_AWCACHE(m_axi_edges_3_AWCACHE),
    .m_axi_AWID(m_axi_edges_3_AWID),
    .m_axi_AWLEN(m_axi_edges_3_AWLEN),
    .m_axi_AWLOCK(m_axi_edges_3_AWLOCK),
    .m_axi_AWPROT(m_axi_edges_3_AWPROT),
    .m_axi_AWQOS(m_axi_edges_3_AWQOS),
    .m_axi_AWREADY(m_axi_edges_3_AWREADY),
    .m_axi_AWREGION(m_axi_edges_3_AWREGION),
    .m_axi_AWSIZE(m_axi_edges_3_AWSIZE),
    .m_axi_AWUSER(m_axi_edges_3_AWUSER),
    .m_axi_AWVALID(m_axi_edges_3_AWVALID),
    .m_axi_BID(m_axi_edges_3_BID),
    .m_axi_BREADY(m_axi_edges_3_BREADY),
    .m_axi_BRESP(m_axi_edges_3_BRESP),
    .m_axi_BUSER(m_axi_edges_3_BUSER),
    .m_axi_BVALID(m_axi_edges_3_BVALID),
    .m_axi_RDATA(m_axi_edges_3_RDATA),
    .m_axi_RID(m_axi_edges_3_RID),
    .m_axi_RLAST(m_axi_edges_3_RLAST),
    .m_axi_RREADY(m_axi_edges_3_RREADY),
    .m_axi_RRESP(m_axi_edges_3_RRESP),
    .m_axi_RUSER(m_axi_edges_3_RUSER),
    .m_axi_RVALID(m_axi_edges_3_RVALID),
    .m_axi_WDATA(m_axi_edges_3_WDATA),
    .m_axi_WID(m_axi_edges_3_WID),
    .m_axi_WLAST(m_axi_edges_3_WLAST),
    .m_axi_WREADY(m_axi_edges_3_WREADY),
    .m_axi_WSTRB(m_axi_edges_3_WSTRB),
    .m_axi_WUSER(m_axi_edges_3_WUSER),
    .m_axi_WVALID(m_axi_edges_3_WVALID),
    .read_addr_din(edges_3__q2 + {edges_3_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(edges_3_read_addr__full_n),
    .read_addr_write(edges_3_read_addr__write),
    .read_data_dout(edges_3_read_data__dout),
    .read_data_empty_n(edges_3_read_data__empty_n),
    .read_data_read(edges_3_read_data__read),
    .write_addr_din('d0),
    .write_addr_full_n(),
    .write_addr_write(1'b0),
    .write_data_din('d0),
    .write_data_full_n(),
    .write_data_write(1'b0)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  edges_4__m_axi
  (
    .clk(ap_clk),
    .rst(edges_4__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_edges_4_ARADDR),
    .m_axi_ARBURST(m_axi_edges_4_ARBURST),
    .m_axi_ARCACHE(m_axi_edges_4_ARCACHE),
    .m_axi_ARID(m_axi_edges_4_ARID),
    .m_axi_ARLEN(m_axi_edges_4_ARLEN),
    .m_axi_ARLOCK(m_axi_edges_4_ARLOCK),
    .m_axi_ARPROT(m_axi_edges_4_ARPROT),
    .m_axi_ARQOS(m_axi_edges_4_ARQOS),
    .m_axi_ARREADY(m_axi_edges_4_ARREADY),
    .m_axi_ARREGION(m_axi_edges_4_ARREGION),
    .m_axi_ARSIZE(m_axi_edges_4_ARSIZE),
    .m_axi_ARUSER(m_axi_edges_4_ARUSER),
    .m_axi_ARVALID(m_axi_edges_4_ARVALID),
    .m_axi_AWADDR(m_axi_edges_4_AWADDR),
    .m_axi_AWBURST(m_axi_edges_4_AWBURST),
    .m_axi_AWCACHE(m_axi_edges_4_AWCACHE),
    .m_axi_AWID(m_axi_edges_4_AWID),
    .m_axi_AWLEN(m_axi_edges_4_AWLEN),
    .m_axi_AWLOCK(m_axi_edges_4_AWLOCK),
    .m_axi_AWPROT(m_axi_edges_4_AWPROT),
    .m_axi_AWQOS(m_axi_edges_4_AWQOS),
    .m_axi_AWREADY(m_axi_edges_4_AWREADY),
    .m_axi_AWREGION(m_axi_edges_4_AWREGION),
    .m_axi_AWSIZE(m_axi_edges_4_AWSIZE),
    .m_axi_AWUSER(m_axi_edges_4_AWUSER),
    .m_axi_AWVALID(m_axi_edges_4_AWVALID),
    .m_axi_BID(m_axi_edges_4_BID),
    .m_axi_BREADY(m_axi_edges_4_BREADY),
    .m_axi_BRESP(m_axi_edges_4_BRESP),
    .m_axi_BUSER(m_axi_edges_4_BUSER),
    .m_axi_BVALID(m_axi_edges_4_BVALID),
    .m_axi_RDATA(m_axi_edges_4_RDATA),
    .m_axi_RID(m_axi_edges_4_RID),
    .m_axi_RLAST(m_axi_edges_4_RLAST),
    .m_axi_RREADY(m_axi_edges_4_RREADY),
    .m_axi_RRESP(m_axi_edges_4_RRESP),
    .m_axi_RUSER(m_axi_edges_4_RUSER),
    .m_axi_RVALID(m_axi_edges_4_RVALID),
    .m_axi_WDATA(m_axi_edges_4_WDATA),
    .m_axi_WID(m_axi_edges_4_WID),
    .m_axi_WLAST(m_axi_edges_4_WLAST),
    .m_axi_WREADY(m_axi_edges_4_WREADY),
    .m_axi_WSTRB(m_axi_edges_4_WSTRB),
    .m_axi_WUSER(m_axi_edges_4_WUSER),
    .m_axi_WVALID(m_axi_edges_4_WVALID),
    .read_addr_din(edges_4__q2 + {edges_4_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(edges_4_read_addr__full_n),
    .read_addr_write(edges_4_read_addr__write),
    .read_data_dout(edges_4_read_data__dout),
    .read_data_empty_n(edges_4_read_data__empty_n),
    .read_data_read(edges_4_read_data__read),
    .write_addr_din('d0),
    .write_addr_full_n(),
    .write_addr_write(1'b0),
    .write_data_din('d0),
    .write_data_full_n(),
    .write_data_write(1'b0)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  edges_5__m_axi
  (
    .clk(ap_clk),
    .rst(edges_5__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_edges_5_ARADDR),
    .m_axi_ARBURST(m_axi_edges_5_ARBURST),
    .m_axi_ARCACHE(m_axi_edges_5_ARCACHE),
    .m_axi_ARID(m_axi_edges_5_ARID),
    .m_axi_ARLEN(m_axi_edges_5_ARLEN),
    .m_axi_ARLOCK(m_axi_edges_5_ARLOCK),
    .m_axi_ARPROT(m_axi_edges_5_ARPROT),
    .m_axi_ARQOS(m_axi_edges_5_ARQOS),
    .m_axi_ARREADY(m_axi_edges_5_ARREADY),
    .m_axi_ARREGION(m_axi_edges_5_ARREGION),
    .m_axi_ARSIZE(m_axi_edges_5_ARSIZE),
    .m_axi_ARUSER(m_axi_edges_5_ARUSER),
    .m_axi_ARVALID(m_axi_edges_5_ARVALID),
    .m_axi_AWADDR(m_axi_edges_5_AWADDR),
    .m_axi_AWBURST(m_axi_edges_5_AWBURST),
    .m_axi_AWCACHE(m_axi_edges_5_AWCACHE),
    .m_axi_AWID(m_axi_edges_5_AWID),
    .m_axi_AWLEN(m_axi_edges_5_AWLEN),
    .m_axi_AWLOCK(m_axi_edges_5_AWLOCK),
    .m_axi_AWPROT(m_axi_edges_5_AWPROT),
    .m_axi_AWQOS(m_axi_edges_5_AWQOS),
    .m_axi_AWREADY(m_axi_edges_5_AWREADY),
    .m_axi_AWREGION(m_axi_edges_5_AWREGION),
    .m_axi_AWSIZE(m_axi_edges_5_AWSIZE),
    .m_axi_AWUSER(m_axi_edges_5_AWUSER),
    .m_axi_AWVALID(m_axi_edges_5_AWVALID),
    .m_axi_BID(m_axi_edges_5_BID),
    .m_axi_BREADY(m_axi_edges_5_BREADY),
    .m_axi_BRESP(m_axi_edges_5_BRESP),
    .m_axi_BUSER(m_axi_edges_5_BUSER),
    .m_axi_BVALID(m_axi_edges_5_BVALID),
    .m_axi_RDATA(m_axi_edges_5_RDATA),
    .m_axi_RID(m_axi_edges_5_RID),
    .m_axi_RLAST(m_axi_edges_5_RLAST),
    .m_axi_RREADY(m_axi_edges_5_RREADY),
    .m_axi_RRESP(m_axi_edges_5_RRESP),
    .m_axi_RUSER(m_axi_edges_5_RUSER),
    .m_axi_RVALID(m_axi_edges_5_RVALID),
    .m_axi_WDATA(m_axi_edges_5_WDATA),
    .m_axi_WID(m_axi_edges_5_WID),
    .m_axi_WLAST(m_axi_edges_5_WLAST),
    .m_axi_WREADY(m_axi_edges_5_WREADY),
    .m_axi_WSTRB(m_axi_edges_5_WSTRB),
    .m_axi_WUSER(m_axi_edges_5_WUSER),
    .m_axi_WVALID(m_axi_edges_5_WVALID),
    .read_addr_din(edges_5__q2 + {edges_5_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(edges_5_read_addr__full_n),
    .read_addr_write(edges_5_read_addr__write),
    .read_data_dout(edges_5_read_data__dout),
    .read_data_empty_n(edges_5_read_data__empty_n),
    .read_data_read(edges_5_read_data__read),
    .write_addr_din('d0),
    .write_addr_full_n(),
    .write_addr_write(1'b0),
    .write_data_din('d0),
    .write_data_full_n(),
    .write_data_write(1'b0)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  edges_6__m_axi
  (
    .clk(ap_clk),
    .rst(edges_6__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_edges_6_ARADDR),
    .m_axi_ARBURST(m_axi_edges_6_ARBURST),
    .m_axi_ARCACHE(m_axi_edges_6_ARCACHE),
    .m_axi_ARID(m_axi_edges_6_ARID),
    .m_axi_ARLEN(m_axi_edges_6_ARLEN),
    .m_axi_ARLOCK(m_axi_edges_6_ARLOCK),
    .m_axi_ARPROT(m_axi_edges_6_ARPROT),
    .m_axi_ARQOS(m_axi_edges_6_ARQOS),
    .m_axi_ARREADY(m_axi_edges_6_ARREADY),
    .m_axi_ARREGION(m_axi_edges_6_ARREGION),
    .m_axi_ARSIZE(m_axi_edges_6_ARSIZE),
    .m_axi_ARUSER(m_axi_edges_6_ARUSER),
    .m_axi_ARVALID(m_axi_edges_6_ARVALID),
    .m_axi_AWADDR(m_axi_edges_6_AWADDR),
    .m_axi_AWBURST(m_axi_edges_6_AWBURST),
    .m_axi_AWCACHE(m_axi_edges_6_AWCACHE),
    .m_axi_AWID(m_axi_edges_6_AWID),
    .m_axi_AWLEN(m_axi_edges_6_AWLEN),
    .m_axi_AWLOCK(m_axi_edges_6_AWLOCK),
    .m_axi_AWPROT(m_axi_edges_6_AWPROT),
    .m_axi_AWQOS(m_axi_edges_6_AWQOS),
    .m_axi_AWREADY(m_axi_edges_6_AWREADY),
    .m_axi_AWREGION(m_axi_edges_6_AWREGION),
    .m_axi_AWSIZE(m_axi_edges_6_AWSIZE),
    .m_axi_AWUSER(m_axi_edges_6_AWUSER),
    .m_axi_AWVALID(m_axi_edges_6_AWVALID),
    .m_axi_BID(m_axi_edges_6_BID),
    .m_axi_BREADY(m_axi_edges_6_BREADY),
    .m_axi_BRESP(m_axi_edges_6_BRESP),
    .m_axi_BUSER(m_axi_edges_6_BUSER),
    .m_axi_BVALID(m_axi_edges_6_BVALID),
    .m_axi_RDATA(m_axi_edges_6_RDATA),
    .m_axi_RID(m_axi_edges_6_RID),
    .m_axi_RLAST(m_axi_edges_6_RLAST),
    .m_axi_RREADY(m_axi_edges_6_RREADY),
    .m_axi_RRESP(m_axi_edges_6_RRESP),
    .m_axi_RUSER(m_axi_edges_6_RUSER),
    .m_axi_RVALID(m_axi_edges_6_RVALID),
    .m_axi_WDATA(m_axi_edges_6_WDATA),
    .m_axi_WID(m_axi_edges_6_WID),
    .m_axi_WLAST(m_axi_edges_6_WLAST),
    .m_axi_WREADY(m_axi_edges_6_WREADY),
    .m_axi_WSTRB(m_axi_edges_6_WSTRB),
    .m_axi_WUSER(m_axi_edges_6_WUSER),
    .m_axi_WVALID(m_axi_edges_6_WVALID),
    .read_addr_din(edges_6__q2 + {edges_6_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(edges_6_read_addr__full_n),
    .read_addr_write(edges_6_read_addr__write),
    .read_data_dout(edges_6_read_data__dout),
    .read_data_empty_n(edges_6_read_data__empty_n),
    .read_data_read(edges_6_read_data__read),
    .write_addr_din('d0),
    .write_addr_full_n(),
    .write_addr_write(1'b0),
    .write_data_din('d0),
    .write_data_full_n(),
    .write_data_write(1'b0)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  edges_7__m_axi
  (
    .clk(ap_clk),
    .rst(edges_7__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_edges_7_ARADDR),
    .m_axi_ARBURST(m_axi_edges_7_ARBURST),
    .m_axi_ARCACHE(m_axi_edges_7_ARCACHE),
    .m_axi_ARID(m_axi_edges_7_ARID),
    .m_axi_ARLEN(m_axi_edges_7_ARLEN),
    .m_axi_ARLOCK(m_axi_edges_7_ARLOCK),
    .m_axi_ARPROT(m_axi_edges_7_ARPROT),
    .m_axi_ARQOS(m_axi_edges_7_ARQOS),
    .m_axi_ARREADY(m_axi_edges_7_ARREADY),
    .m_axi_ARREGION(m_axi_edges_7_ARREGION),
    .m_axi_ARSIZE(m_axi_edges_7_ARSIZE),
    .m_axi_ARUSER(m_axi_edges_7_ARUSER),
    .m_axi_ARVALID(m_axi_edges_7_ARVALID),
    .m_axi_AWADDR(m_axi_edges_7_AWADDR),
    .m_axi_AWBURST(m_axi_edges_7_AWBURST),
    .m_axi_AWCACHE(m_axi_edges_7_AWCACHE),
    .m_axi_AWID(m_axi_edges_7_AWID),
    .m_axi_AWLEN(m_axi_edges_7_AWLEN),
    .m_axi_AWLOCK(m_axi_edges_7_AWLOCK),
    .m_axi_AWPROT(m_axi_edges_7_AWPROT),
    .m_axi_AWQOS(m_axi_edges_7_AWQOS),
    .m_axi_AWREADY(m_axi_edges_7_AWREADY),
    .m_axi_AWREGION(m_axi_edges_7_AWREGION),
    .m_axi_AWSIZE(m_axi_edges_7_AWSIZE),
    .m_axi_AWUSER(m_axi_edges_7_AWUSER),
    .m_axi_AWVALID(m_axi_edges_7_AWVALID),
    .m_axi_BID(m_axi_edges_7_BID),
    .m_axi_BREADY(m_axi_edges_7_BREADY),
    .m_axi_BRESP(m_axi_edges_7_BRESP),
    .m_axi_BUSER(m_axi_edges_7_BUSER),
    .m_axi_BVALID(m_axi_edges_7_BVALID),
    .m_axi_RDATA(m_axi_edges_7_RDATA),
    .m_axi_RID(m_axi_edges_7_RID),
    .m_axi_RLAST(m_axi_edges_7_RLAST),
    .m_axi_RREADY(m_axi_edges_7_RREADY),
    .m_axi_RRESP(m_axi_edges_7_RRESP),
    .m_axi_RUSER(m_axi_edges_7_RUSER),
    .m_axi_RVALID(m_axi_edges_7_RVALID),
    .m_axi_WDATA(m_axi_edges_7_WDATA),
    .m_axi_WID(m_axi_edges_7_WID),
    .m_axi_WLAST(m_axi_edges_7_WLAST),
    .m_axi_WREADY(m_axi_edges_7_WREADY),
    .m_axi_WSTRB(m_axi_edges_7_WSTRB),
    .m_axi_WUSER(m_axi_edges_7_WUSER),
    .m_axi_WVALID(m_axi_edges_7_WVALID),
    .read_addr_din(edges_7__q2 + {edges_7_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(edges_7_read_addr__full_n),
    .read_addr_write(edges_7_read_addr__write),
    .read_data_dout(edges_7_read_data__dout),
    .read_data_empty_n(edges_7_read_data__empty_n),
    .read_data_read(edges_7_read_data__read),
    .write_addr_din('d0),
    .write_addr_full_n(),
    .write_addr_write(1'b0),
    .write_data_din('d0),
    .write_data_full_n(),
    .write_data_write(1'b0)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  updates_0__m_axi
  (
    .clk(ap_clk),
    .rst(updates_0__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_updates_0_ARADDR),
    .m_axi_ARBURST(m_axi_updates_0_ARBURST),
    .m_axi_ARCACHE(m_axi_updates_0_ARCACHE),
    .m_axi_ARID(m_axi_updates_0_ARID),
    .m_axi_ARLEN(m_axi_updates_0_ARLEN),
    .m_axi_ARLOCK(m_axi_updates_0_ARLOCK),
    .m_axi_ARPROT(m_axi_updates_0_ARPROT),
    .m_axi_ARQOS(m_axi_updates_0_ARQOS),
    .m_axi_ARREADY(m_axi_updates_0_ARREADY),
    .m_axi_ARREGION(m_axi_updates_0_ARREGION),
    .m_axi_ARSIZE(m_axi_updates_0_ARSIZE),
    .m_axi_ARUSER(m_axi_updates_0_ARUSER),
    .m_axi_ARVALID(m_axi_updates_0_ARVALID),
    .m_axi_AWADDR(m_axi_updates_0_AWADDR),
    .m_axi_AWBURST(m_axi_updates_0_AWBURST),
    .m_axi_AWCACHE(m_axi_updates_0_AWCACHE),
    .m_axi_AWID(m_axi_updates_0_AWID),
    .m_axi_AWLEN(m_axi_updates_0_AWLEN),
    .m_axi_AWLOCK(m_axi_updates_0_AWLOCK),
    .m_axi_AWPROT(m_axi_updates_0_AWPROT),
    .m_axi_AWQOS(m_axi_updates_0_AWQOS),
    .m_axi_AWREADY(m_axi_updates_0_AWREADY),
    .m_axi_AWREGION(m_axi_updates_0_AWREGION),
    .m_axi_AWSIZE(m_axi_updates_0_AWSIZE),
    .m_axi_AWUSER(m_axi_updates_0_AWUSER),
    .m_axi_AWVALID(m_axi_updates_0_AWVALID),
    .m_axi_BID(m_axi_updates_0_BID),
    .m_axi_BREADY(m_axi_updates_0_BREADY),
    .m_axi_BRESP(m_axi_updates_0_BRESP),
    .m_axi_BUSER(m_axi_updates_0_BUSER),
    .m_axi_BVALID(m_axi_updates_0_BVALID),
    .m_axi_RDATA(m_axi_updates_0_RDATA),
    .m_axi_RID(m_axi_updates_0_RID),
    .m_axi_RLAST(m_axi_updates_0_RLAST),
    .m_axi_RREADY(m_axi_updates_0_RREADY),
    .m_axi_RRESP(m_axi_updates_0_RRESP),
    .m_axi_RUSER(m_axi_updates_0_RUSER),
    .m_axi_RVALID(m_axi_updates_0_RVALID),
    .m_axi_WDATA(m_axi_updates_0_WDATA),
    .m_axi_WID(m_axi_updates_0_WID),
    .m_axi_WLAST(m_axi_updates_0_WLAST),
    .m_axi_WREADY(m_axi_updates_0_WREADY),
    .m_axi_WSTRB(m_axi_updates_0_WSTRB),
    .m_axi_WUSER(m_axi_updates_0_WUSER),
    .m_axi_WVALID(m_axi_updates_0_WVALID),
    .read_addr_din(updates_0__q2 + {updates_0_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(updates_0_read_addr__full_n),
    .read_addr_write(updates_0_read_addr__write),
    .read_data_dout(updates_0_read_data__dout),
    .read_data_empty_n(updates_0_read_data__empty_n),
    .read_data_read(updates_0_read_data__read),
    .write_addr_din(updates_0__q2 + {updates_0_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(updates_0_write_addr__full_n),
    .write_addr_write(updates_0_write_addr__write),
    .write_data_din(updates_0_write_data__din),
    .write_data_full_n(updates_0_write_data__full_n),
    .write_data_write(updates_0_write_data__write)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  updates_1__m_axi
  (
    .clk(ap_clk),
    .rst(updates_1__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_updates_1_ARADDR),
    .m_axi_ARBURST(m_axi_updates_1_ARBURST),
    .m_axi_ARCACHE(m_axi_updates_1_ARCACHE),
    .m_axi_ARID(m_axi_updates_1_ARID),
    .m_axi_ARLEN(m_axi_updates_1_ARLEN),
    .m_axi_ARLOCK(m_axi_updates_1_ARLOCK),
    .m_axi_ARPROT(m_axi_updates_1_ARPROT),
    .m_axi_ARQOS(m_axi_updates_1_ARQOS),
    .m_axi_ARREADY(m_axi_updates_1_ARREADY),
    .m_axi_ARREGION(m_axi_updates_1_ARREGION),
    .m_axi_ARSIZE(m_axi_updates_1_ARSIZE),
    .m_axi_ARUSER(m_axi_updates_1_ARUSER),
    .m_axi_ARVALID(m_axi_updates_1_ARVALID),
    .m_axi_AWADDR(m_axi_updates_1_AWADDR),
    .m_axi_AWBURST(m_axi_updates_1_AWBURST),
    .m_axi_AWCACHE(m_axi_updates_1_AWCACHE),
    .m_axi_AWID(m_axi_updates_1_AWID),
    .m_axi_AWLEN(m_axi_updates_1_AWLEN),
    .m_axi_AWLOCK(m_axi_updates_1_AWLOCK),
    .m_axi_AWPROT(m_axi_updates_1_AWPROT),
    .m_axi_AWQOS(m_axi_updates_1_AWQOS),
    .m_axi_AWREADY(m_axi_updates_1_AWREADY),
    .m_axi_AWREGION(m_axi_updates_1_AWREGION),
    .m_axi_AWSIZE(m_axi_updates_1_AWSIZE),
    .m_axi_AWUSER(m_axi_updates_1_AWUSER),
    .m_axi_AWVALID(m_axi_updates_1_AWVALID),
    .m_axi_BID(m_axi_updates_1_BID),
    .m_axi_BREADY(m_axi_updates_1_BREADY),
    .m_axi_BRESP(m_axi_updates_1_BRESP),
    .m_axi_BUSER(m_axi_updates_1_BUSER),
    .m_axi_BVALID(m_axi_updates_1_BVALID),
    .m_axi_RDATA(m_axi_updates_1_RDATA),
    .m_axi_RID(m_axi_updates_1_RID),
    .m_axi_RLAST(m_axi_updates_1_RLAST),
    .m_axi_RREADY(m_axi_updates_1_RREADY),
    .m_axi_RRESP(m_axi_updates_1_RRESP),
    .m_axi_RUSER(m_axi_updates_1_RUSER),
    .m_axi_RVALID(m_axi_updates_1_RVALID),
    .m_axi_WDATA(m_axi_updates_1_WDATA),
    .m_axi_WID(m_axi_updates_1_WID),
    .m_axi_WLAST(m_axi_updates_1_WLAST),
    .m_axi_WREADY(m_axi_updates_1_WREADY),
    .m_axi_WSTRB(m_axi_updates_1_WSTRB),
    .m_axi_WUSER(m_axi_updates_1_WUSER),
    .m_axi_WVALID(m_axi_updates_1_WVALID),
    .read_addr_din(updates_1__q2 + {updates_1_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(updates_1_read_addr__full_n),
    .read_addr_write(updates_1_read_addr__write),
    .read_data_dout(updates_1_read_data__dout),
    .read_data_empty_n(updates_1_read_data__empty_n),
    .read_data_read(updates_1_read_data__read),
    .write_addr_din(updates_1__q2 + {updates_1_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(updates_1_write_addr__full_n),
    .write_addr_write(updates_1_write_addr__write),
    .write_data_din(updates_1_write_data__din),
    .write_data_full_n(updates_1_write_data__full_n),
    .write_data_write(updates_1_write_data__write)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  updates_2__m_axi
  (
    .clk(ap_clk),
    .rst(updates_2__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_updates_2_ARADDR),
    .m_axi_ARBURST(m_axi_updates_2_ARBURST),
    .m_axi_ARCACHE(m_axi_updates_2_ARCACHE),
    .m_axi_ARID(m_axi_updates_2_ARID),
    .m_axi_ARLEN(m_axi_updates_2_ARLEN),
    .m_axi_ARLOCK(m_axi_updates_2_ARLOCK),
    .m_axi_ARPROT(m_axi_updates_2_ARPROT),
    .m_axi_ARQOS(m_axi_updates_2_ARQOS),
    .m_axi_ARREADY(m_axi_updates_2_ARREADY),
    .m_axi_ARREGION(m_axi_updates_2_ARREGION),
    .m_axi_ARSIZE(m_axi_updates_2_ARSIZE),
    .m_axi_ARUSER(m_axi_updates_2_ARUSER),
    .m_axi_ARVALID(m_axi_updates_2_ARVALID),
    .m_axi_AWADDR(m_axi_updates_2_AWADDR),
    .m_axi_AWBURST(m_axi_updates_2_AWBURST),
    .m_axi_AWCACHE(m_axi_updates_2_AWCACHE),
    .m_axi_AWID(m_axi_updates_2_AWID),
    .m_axi_AWLEN(m_axi_updates_2_AWLEN),
    .m_axi_AWLOCK(m_axi_updates_2_AWLOCK),
    .m_axi_AWPROT(m_axi_updates_2_AWPROT),
    .m_axi_AWQOS(m_axi_updates_2_AWQOS),
    .m_axi_AWREADY(m_axi_updates_2_AWREADY),
    .m_axi_AWREGION(m_axi_updates_2_AWREGION),
    .m_axi_AWSIZE(m_axi_updates_2_AWSIZE),
    .m_axi_AWUSER(m_axi_updates_2_AWUSER),
    .m_axi_AWVALID(m_axi_updates_2_AWVALID),
    .m_axi_BID(m_axi_updates_2_BID),
    .m_axi_BREADY(m_axi_updates_2_BREADY),
    .m_axi_BRESP(m_axi_updates_2_BRESP),
    .m_axi_BUSER(m_axi_updates_2_BUSER),
    .m_axi_BVALID(m_axi_updates_2_BVALID),
    .m_axi_RDATA(m_axi_updates_2_RDATA),
    .m_axi_RID(m_axi_updates_2_RID),
    .m_axi_RLAST(m_axi_updates_2_RLAST),
    .m_axi_RREADY(m_axi_updates_2_RREADY),
    .m_axi_RRESP(m_axi_updates_2_RRESP),
    .m_axi_RUSER(m_axi_updates_2_RUSER),
    .m_axi_RVALID(m_axi_updates_2_RVALID),
    .m_axi_WDATA(m_axi_updates_2_WDATA),
    .m_axi_WID(m_axi_updates_2_WID),
    .m_axi_WLAST(m_axi_updates_2_WLAST),
    .m_axi_WREADY(m_axi_updates_2_WREADY),
    .m_axi_WSTRB(m_axi_updates_2_WSTRB),
    .m_axi_WUSER(m_axi_updates_2_WUSER),
    .m_axi_WVALID(m_axi_updates_2_WVALID),
    .read_addr_din(updates_2__q2 + {updates_2_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(updates_2_read_addr__full_n),
    .read_addr_write(updates_2_read_addr__write),
    .read_data_dout(updates_2_read_data__dout),
    .read_data_empty_n(updates_2_read_data__empty_n),
    .read_data_read(updates_2_read_data__read),
    .write_addr_din(updates_2__q2 + {updates_2_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(updates_2_write_addr__full_n),
    .write_addr_write(updates_2_write_addr__write),
    .write_data_din(updates_2_write_data__din),
    .write_data_full_n(updates_2_write_data__full_n),
    .write_data_write(updates_2_write_data__write)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  updates_3__m_axi
  (
    .clk(ap_clk),
    .rst(updates_3__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_updates_3_ARADDR),
    .m_axi_ARBURST(m_axi_updates_3_ARBURST),
    .m_axi_ARCACHE(m_axi_updates_3_ARCACHE),
    .m_axi_ARID(m_axi_updates_3_ARID),
    .m_axi_ARLEN(m_axi_updates_3_ARLEN),
    .m_axi_ARLOCK(m_axi_updates_3_ARLOCK),
    .m_axi_ARPROT(m_axi_updates_3_ARPROT),
    .m_axi_ARQOS(m_axi_updates_3_ARQOS),
    .m_axi_ARREADY(m_axi_updates_3_ARREADY),
    .m_axi_ARREGION(m_axi_updates_3_ARREGION),
    .m_axi_ARSIZE(m_axi_updates_3_ARSIZE),
    .m_axi_ARUSER(m_axi_updates_3_ARUSER),
    .m_axi_ARVALID(m_axi_updates_3_ARVALID),
    .m_axi_AWADDR(m_axi_updates_3_AWADDR),
    .m_axi_AWBURST(m_axi_updates_3_AWBURST),
    .m_axi_AWCACHE(m_axi_updates_3_AWCACHE),
    .m_axi_AWID(m_axi_updates_3_AWID),
    .m_axi_AWLEN(m_axi_updates_3_AWLEN),
    .m_axi_AWLOCK(m_axi_updates_3_AWLOCK),
    .m_axi_AWPROT(m_axi_updates_3_AWPROT),
    .m_axi_AWQOS(m_axi_updates_3_AWQOS),
    .m_axi_AWREADY(m_axi_updates_3_AWREADY),
    .m_axi_AWREGION(m_axi_updates_3_AWREGION),
    .m_axi_AWSIZE(m_axi_updates_3_AWSIZE),
    .m_axi_AWUSER(m_axi_updates_3_AWUSER),
    .m_axi_AWVALID(m_axi_updates_3_AWVALID),
    .m_axi_BID(m_axi_updates_3_BID),
    .m_axi_BREADY(m_axi_updates_3_BREADY),
    .m_axi_BRESP(m_axi_updates_3_BRESP),
    .m_axi_BUSER(m_axi_updates_3_BUSER),
    .m_axi_BVALID(m_axi_updates_3_BVALID),
    .m_axi_RDATA(m_axi_updates_3_RDATA),
    .m_axi_RID(m_axi_updates_3_RID),
    .m_axi_RLAST(m_axi_updates_3_RLAST),
    .m_axi_RREADY(m_axi_updates_3_RREADY),
    .m_axi_RRESP(m_axi_updates_3_RRESP),
    .m_axi_RUSER(m_axi_updates_3_RUSER),
    .m_axi_RVALID(m_axi_updates_3_RVALID),
    .m_axi_WDATA(m_axi_updates_3_WDATA),
    .m_axi_WID(m_axi_updates_3_WID),
    .m_axi_WLAST(m_axi_updates_3_WLAST),
    .m_axi_WREADY(m_axi_updates_3_WREADY),
    .m_axi_WSTRB(m_axi_updates_3_WSTRB),
    .m_axi_WUSER(m_axi_updates_3_WUSER),
    .m_axi_WVALID(m_axi_updates_3_WVALID),
    .read_addr_din(updates_3__q2 + {updates_3_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(updates_3_read_addr__full_n),
    .read_addr_write(updates_3_read_addr__write),
    .read_data_dout(updates_3_read_data__dout),
    .read_data_empty_n(updates_3_read_data__empty_n),
    .read_data_read(updates_3_read_data__read),
    .write_addr_din(updates_3__q2 + {updates_3_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(updates_3_write_addr__full_n),
    .write_addr_write(updates_3_write_addr__write),
    .write_data_din(updates_3_write_data__din),
    .write_data_full_n(updates_3_write_data__full_n),
    .write_data_write(updates_3_write_data__write)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  updates_4__m_axi
  (
    .clk(ap_clk),
    .rst(updates_4__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_updates_4_ARADDR),
    .m_axi_ARBURST(m_axi_updates_4_ARBURST),
    .m_axi_ARCACHE(m_axi_updates_4_ARCACHE),
    .m_axi_ARID(m_axi_updates_4_ARID),
    .m_axi_ARLEN(m_axi_updates_4_ARLEN),
    .m_axi_ARLOCK(m_axi_updates_4_ARLOCK),
    .m_axi_ARPROT(m_axi_updates_4_ARPROT),
    .m_axi_ARQOS(m_axi_updates_4_ARQOS),
    .m_axi_ARREADY(m_axi_updates_4_ARREADY),
    .m_axi_ARREGION(m_axi_updates_4_ARREGION),
    .m_axi_ARSIZE(m_axi_updates_4_ARSIZE),
    .m_axi_ARUSER(m_axi_updates_4_ARUSER),
    .m_axi_ARVALID(m_axi_updates_4_ARVALID),
    .m_axi_AWADDR(m_axi_updates_4_AWADDR),
    .m_axi_AWBURST(m_axi_updates_4_AWBURST),
    .m_axi_AWCACHE(m_axi_updates_4_AWCACHE),
    .m_axi_AWID(m_axi_updates_4_AWID),
    .m_axi_AWLEN(m_axi_updates_4_AWLEN),
    .m_axi_AWLOCK(m_axi_updates_4_AWLOCK),
    .m_axi_AWPROT(m_axi_updates_4_AWPROT),
    .m_axi_AWQOS(m_axi_updates_4_AWQOS),
    .m_axi_AWREADY(m_axi_updates_4_AWREADY),
    .m_axi_AWREGION(m_axi_updates_4_AWREGION),
    .m_axi_AWSIZE(m_axi_updates_4_AWSIZE),
    .m_axi_AWUSER(m_axi_updates_4_AWUSER),
    .m_axi_AWVALID(m_axi_updates_4_AWVALID),
    .m_axi_BID(m_axi_updates_4_BID),
    .m_axi_BREADY(m_axi_updates_4_BREADY),
    .m_axi_BRESP(m_axi_updates_4_BRESP),
    .m_axi_BUSER(m_axi_updates_4_BUSER),
    .m_axi_BVALID(m_axi_updates_4_BVALID),
    .m_axi_RDATA(m_axi_updates_4_RDATA),
    .m_axi_RID(m_axi_updates_4_RID),
    .m_axi_RLAST(m_axi_updates_4_RLAST),
    .m_axi_RREADY(m_axi_updates_4_RREADY),
    .m_axi_RRESP(m_axi_updates_4_RRESP),
    .m_axi_RUSER(m_axi_updates_4_RUSER),
    .m_axi_RVALID(m_axi_updates_4_RVALID),
    .m_axi_WDATA(m_axi_updates_4_WDATA),
    .m_axi_WID(m_axi_updates_4_WID),
    .m_axi_WLAST(m_axi_updates_4_WLAST),
    .m_axi_WREADY(m_axi_updates_4_WREADY),
    .m_axi_WSTRB(m_axi_updates_4_WSTRB),
    .m_axi_WUSER(m_axi_updates_4_WUSER),
    .m_axi_WVALID(m_axi_updates_4_WVALID),
    .read_addr_din(updates_4__q2 + {updates_4_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(updates_4_read_addr__full_n),
    .read_addr_write(updates_4_read_addr__write),
    .read_data_dout(updates_4_read_data__dout),
    .read_data_empty_n(updates_4_read_data__empty_n),
    .read_data_read(updates_4_read_data__read),
    .write_addr_din(updates_4__q2 + {updates_4_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(updates_4_write_addr__full_n),
    .write_addr_write(updates_4_write_addr__write),
    .write_data_din(updates_4_write_data__din),
    .write_data_full_n(updates_4_write_data__full_n),
    .write_data_write(updates_4_write_data__write)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  updates_5__m_axi
  (
    .clk(ap_clk),
    .rst(updates_5__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_updates_5_ARADDR),
    .m_axi_ARBURST(m_axi_updates_5_ARBURST),
    .m_axi_ARCACHE(m_axi_updates_5_ARCACHE),
    .m_axi_ARID(m_axi_updates_5_ARID),
    .m_axi_ARLEN(m_axi_updates_5_ARLEN),
    .m_axi_ARLOCK(m_axi_updates_5_ARLOCK),
    .m_axi_ARPROT(m_axi_updates_5_ARPROT),
    .m_axi_ARQOS(m_axi_updates_5_ARQOS),
    .m_axi_ARREADY(m_axi_updates_5_ARREADY),
    .m_axi_ARREGION(m_axi_updates_5_ARREGION),
    .m_axi_ARSIZE(m_axi_updates_5_ARSIZE),
    .m_axi_ARUSER(m_axi_updates_5_ARUSER),
    .m_axi_ARVALID(m_axi_updates_5_ARVALID),
    .m_axi_AWADDR(m_axi_updates_5_AWADDR),
    .m_axi_AWBURST(m_axi_updates_5_AWBURST),
    .m_axi_AWCACHE(m_axi_updates_5_AWCACHE),
    .m_axi_AWID(m_axi_updates_5_AWID),
    .m_axi_AWLEN(m_axi_updates_5_AWLEN),
    .m_axi_AWLOCK(m_axi_updates_5_AWLOCK),
    .m_axi_AWPROT(m_axi_updates_5_AWPROT),
    .m_axi_AWQOS(m_axi_updates_5_AWQOS),
    .m_axi_AWREADY(m_axi_updates_5_AWREADY),
    .m_axi_AWREGION(m_axi_updates_5_AWREGION),
    .m_axi_AWSIZE(m_axi_updates_5_AWSIZE),
    .m_axi_AWUSER(m_axi_updates_5_AWUSER),
    .m_axi_AWVALID(m_axi_updates_5_AWVALID),
    .m_axi_BID(m_axi_updates_5_BID),
    .m_axi_BREADY(m_axi_updates_5_BREADY),
    .m_axi_BRESP(m_axi_updates_5_BRESP),
    .m_axi_BUSER(m_axi_updates_5_BUSER),
    .m_axi_BVALID(m_axi_updates_5_BVALID),
    .m_axi_RDATA(m_axi_updates_5_RDATA),
    .m_axi_RID(m_axi_updates_5_RID),
    .m_axi_RLAST(m_axi_updates_5_RLAST),
    .m_axi_RREADY(m_axi_updates_5_RREADY),
    .m_axi_RRESP(m_axi_updates_5_RRESP),
    .m_axi_RUSER(m_axi_updates_5_RUSER),
    .m_axi_RVALID(m_axi_updates_5_RVALID),
    .m_axi_WDATA(m_axi_updates_5_WDATA),
    .m_axi_WID(m_axi_updates_5_WID),
    .m_axi_WLAST(m_axi_updates_5_WLAST),
    .m_axi_WREADY(m_axi_updates_5_WREADY),
    .m_axi_WSTRB(m_axi_updates_5_WSTRB),
    .m_axi_WUSER(m_axi_updates_5_WUSER),
    .m_axi_WVALID(m_axi_updates_5_WVALID),
    .read_addr_din(updates_5__q2 + {updates_5_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(updates_5_read_addr__full_n),
    .read_addr_write(updates_5_read_addr__write),
    .read_data_dout(updates_5_read_data__dout),
    .read_data_empty_n(updates_5_read_data__empty_n),
    .read_data_read(updates_5_read_data__read),
    .write_addr_din(updates_5__q2 + {updates_5_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(updates_5_write_addr__full_n),
    .write_addr_write(updates_5_write_addr__write),
    .write_data_din(updates_5_write_data__din),
    .write_data_full_n(updates_5_write_data__full_n),
    .write_data_write(updates_5_write_data__write)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  updates_6__m_axi
  (
    .clk(ap_clk),
    .rst(updates_6__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_updates_6_ARADDR),
    .m_axi_ARBURST(m_axi_updates_6_ARBURST),
    .m_axi_ARCACHE(m_axi_updates_6_ARCACHE),
    .m_axi_ARID(m_axi_updates_6_ARID),
    .m_axi_ARLEN(m_axi_updates_6_ARLEN),
    .m_axi_ARLOCK(m_axi_updates_6_ARLOCK),
    .m_axi_ARPROT(m_axi_updates_6_ARPROT),
    .m_axi_ARQOS(m_axi_updates_6_ARQOS),
    .m_axi_ARREADY(m_axi_updates_6_ARREADY),
    .m_axi_ARREGION(m_axi_updates_6_ARREGION),
    .m_axi_ARSIZE(m_axi_updates_6_ARSIZE),
    .m_axi_ARUSER(m_axi_updates_6_ARUSER),
    .m_axi_ARVALID(m_axi_updates_6_ARVALID),
    .m_axi_AWADDR(m_axi_updates_6_AWADDR),
    .m_axi_AWBURST(m_axi_updates_6_AWBURST),
    .m_axi_AWCACHE(m_axi_updates_6_AWCACHE),
    .m_axi_AWID(m_axi_updates_6_AWID),
    .m_axi_AWLEN(m_axi_updates_6_AWLEN),
    .m_axi_AWLOCK(m_axi_updates_6_AWLOCK),
    .m_axi_AWPROT(m_axi_updates_6_AWPROT),
    .m_axi_AWQOS(m_axi_updates_6_AWQOS),
    .m_axi_AWREADY(m_axi_updates_6_AWREADY),
    .m_axi_AWREGION(m_axi_updates_6_AWREGION),
    .m_axi_AWSIZE(m_axi_updates_6_AWSIZE),
    .m_axi_AWUSER(m_axi_updates_6_AWUSER),
    .m_axi_AWVALID(m_axi_updates_6_AWVALID),
    .m_axi_BID(m_axi_updates_6_BID),
    .m_axi_BREADY(m_axi_updates_6_BREADY),
    .m_axi_BRESP(m_axi_updates_6_BRESP),
    .m_axi_BUSER(m_axi_updates_6_BUSER),
    .m_axi_BVALID(m_axi_updates_6_BVALID),
    .m_axi_RDATA(m_axi_updates_6_RDATA),
    .m_axi_RID(m_axi_updates_6_RID),
    .m_axi_RLAST(m_axi_updates_6_RLAST),
    .m_axi_RREADY(m_axi_updates_6_RREADY),
    .m_axi_RRESP(m_axi_updates_6_RRESP),
    .m_axi_RUSER(m_axi_updates_6_RUSER),
    .m_axi_RVALID(m_axi_updates_6_RVALID),
    .m_axi_WDATA(m_axi_updates_6_WDATA),
    .m_axi_WID(m_axi_updates_6_WID),
    .m_axi_WLAST(m_axi_updates_6_WLAST),
    .m_axi_WREADY(m_axi_updates_6_WREADY),
    .m_axi_WSTRB(m_axi_updates_6_WSTRB),
    .m_axi_WUSER(m_axi_updates_6_WUSER),
    .m_axi_WVALID(m_axi_updates_6_WVALID),
    .read_addr_din(updates_6__q2 + {updates_6_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(updates_6_read_addr__full_n),
    .read_addr_write(updates_6_read_addr__write),
    .read_data_dout(updates_6_read_data__dout),
    .read_data_empty_n(updates_6_read_data__empty_n),
    .read_data_read(updates_6_read_data__read),
    .write_addr_din(updates_6__q2 + {updates_6_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(updates_6_write_addr__full_n),
    .write_addr_write(updates_6_write_addr__write),
    .write_data_din(updates_6_write_data__din),
    .write_data_full_n(updates_6_write_data__full_n),
    .write_data_write(updates_6_write_data__write)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  updates_7__m_axi
  (
    .clk(ap_clk),
    .rst(updates_7__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_updates_7_ARADDR),
    .m_axi_ARBURST(m_axi_updates_7_ARBURST),
    .m_axi_ARCACHE(m_axi_updates_7_ARCACHE),
    .m_axi_ARID(m_axi_updates_7_ARID),
    .m_axi_ARLEN(m_axi_updates_7_ARLEN),
    .m_axi_ARLOCK(m_axi_updates_7_ARLOCK),
    .m_axi_ARPROT(m_axi_updates_7_ARPROT),
    .m_axi_ARQOS(m_axi_updates_7_ARQOS),
    .m_axi_ARREADY(m_axi_updates_7_ARREADY),
    .m_axi_ARREGION(m_axi_updates_7_ARREGION),
    .m_axi_ARSIZE(m_axi_updates_7_ARSIZE),
    .m_axi_ARUSER(m_axi_updates_7_ARUSER),
    .m_axi_ARVALID(m_axi_updates_7_ARVALID),
    .m_axi_AWADDR(m_axi_updates_7_AWADDR),
    .m_axi_AWBURST(m_axi_updates_7_AWBURST),
    .m_axi_AWCACHE(m_axi_updates_7_AWCACHE),
    .m_axi_AWID(m_axi_updates_7_AWID),
    .m_axi_AWLEN(m_axi_updates_7_AWLEN),
    .m_axi_AWLOCK(m_axi_updates_7_AWLOCK),
    .m_axi_AWPROT(m_axi_updates_7_AWPROT),
    .m_axi_AWQOS(m_axi_updates_7_AWQOS),
    .m_axi_AWREADY(m_axi_updates_7_AWREADY),
    .m_axi_AWREGION(m_axi_updates_7_AWREGION),
    .m_axi_AWSIZE(m_axi_updates_7_AWSIZE),
    .m_axi_AWUSER(m_axi_updates_7_AWUSER),
    .m_axi_AWVALID(m_axi_updates_7_AWVALID),
    .m_axi_BID(m_axi_updates_7_BID),
    .m_axi_BREADY(m_axi_updates_7_BREADY),
    .m_axi_BRESP(m_axi_updates_7_BRESP),
    .m_axi_BUSER(m_axi_updates_7_BUSER),
    .m_axi_BVALID(m_axi_updates_7_BVALID),
    .m_axi_RDATA(m_axi_updates_7_RDATA),
    .m_axi_RID(m_axi_updates_7_RID),
    .m_axi_RLAST(m_axi_updates_7_RLAST),
    .m_axi_RREADY(m_axi_updates_7_RREADY),
    .m_axi_RRESP(m_axi_updates_7_RRESP),
    .m_axi_RUSER(m_axi_updates_7_RUSER),
    .m_axi_RVALID(m_axi_updates_7_RVALID),
    .m_axi_WDATA(m_axi_updates_7_WDATA),
    .m_axi_WID(m_axi_updates_7_WID),
    .m_axi_WLAST(m_axi_updates_7_WLAST),
    .m_axi_WREADY(m_axi_updates_7_WREADY),
    .m_axi_WSTRB(m_axi_updates_7_WSTRB),
    .m_axi_WUSER(m_axi_updates_7_WUSER),
    .m_axi_WVALID(m_axi_updates_7_WVALID),
    .read_addr_din(updates_7__q2 + {updates_7_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(updates_7_read_addr__full_n),
    .read_addr_write(updates_7_read_addr__write),
    .read_data_dout(updates_7_read_data__dout),
    .read_data_empty_n(updates_7_read_data__empty_n),
    .read_data_read(updates_7_read_data__read),
    .write_addr_din(updates_7__q2 + {updates_7_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(updates_7_write_addr__full_n),
    .write_addr_write(updates_7_write_addr__write),
    .write_data_din(updates_7_write_data__din),
    .write_data_full_n(updates_7_write_data__full_n),
    .write_data_write(updates_7_write_data__write)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  degrees__m_axi
  (
    .clk(ap_clk),
    .rst(degrees__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_degrees_ARADDR),
    .m_axi_ARBURST(m_axi_degrees_ARBURST),
    .m_axi_ARCACHE(m_axi_degrees_ARCACHE),
    .m_axi_ARID(m_axi_degrees_ARID),
    .m_axi_ARLEN(m_axi_degrees_ARLEN),
    .m_axi_ARLOCK(m_axi_degrees_ARLOCK),
    .m_axi_ARPROT(m_axi_degrees_ARPROT),
    .m_axi_ARQOS(m_axi_degrees_ARQOS),
    .m_axi_ARREADY(m_axi_degrees_ARREADY),
    .m_axi_ARREGION(m_axi_degrees_ARREGION),
    .m_axi_ARSIZE(m_axi_degrees_ARSIZE),
    .m_axi_ARUSER(m_axi_degrees_ARUSER),
    .m_axi_ARVALID(m_axi_degrees_ARVALID),
    .m_axi_AWADDR(m_axi_degrees_AWADDR),
    .m_axi_AWBURST(m_axi_degrees_AWBURST),
    .m_axi_AWCACHE(m_axi_degrees_AWCACHE),
    .m_axi_AWID(m_axi_degrees_AWID),
    .m_axi_AWLEN(m_axi_degrees_AWLEN),
    .m_axi_AWLOCK(m_axi_degrees_AWLOCK),
    .m_axi_AWPROT(m_axi_degrees_AWPROT),
    .m_axi_AWQOS(m_axi_degrees_AWQOS),
    .m_axi_AWREADY(m_axi_degrees_AWREADY),
    .m_axi_AWREGION(m_axi_degrees_AWREGION),
    .m_axi_AWSIZE(m_axi_degrees_AWSIZE),
    .m_axi_AWUSER(m_axi_degrees_AWUSER),
    .m_axi_AWVALID(m_axi_degrees_AWVALID),
    .m_axi_BID(m_axi_degrees_BID),
    .m_axi_BREADY(m_axi_degrees_BREADY),
    .m_axi_BRESP(m_axi_degrees_BRESP),
    .m_axi_BUSER(m_axi_degrees_BUSER),
    .m_axi_BVALID(m_axi_degrees_BVALID),
    .m_axi_RDATA(m_axi_degrees_RDATA),
    .m_axi_RID(m_axi_degrees_RID),
    .m_axi_RLAST(m_axi_degrees_RLAST),
    .m_axi_RREADY(m_axi_degrees_RREADY),
    .m_axi_RRESP(m_axi_degrees_RRESP),
    .m_axi_RUSER(m_axi_degrees_RUSER),
    .m_axi_RVALID(m_axi_degrees_RVALID),
    .m_axi_WDATA(m_axi_degrees_WDATA),
    .m_axi_WID(m_axi_degrees_WID),
    .m_axi_WLAST(m_axi_degrees_WLAST),
    .m_axi_WREADY(m_axi_degrees_WREADY),
    .m_axi_WSTRB(m_axi_degrees_WSTRB),
    .m_axi_WUSER(m_axi_degrees_WUSER),
    .m_axi_WVALID(m_axi_degrees_WVALID),
    .read_addr_din(degrees__q2 + {degrees_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(degrees_read_addr__full_n),
    .read_addr_write(degrees_read_addr__write),
    .read_data_dout(degrees_read_data__dout),
    .read_data_empty_n(degrees_read_data__empty_n),
    .read_data_read(degrees_read_data__read),
    .write_addr_din('d0),
    .write_addr_full_n(),
    .write_addr_write(1'b0),
    .write_data_din('d0),
    .write_data_full_n(),
    .write_data_write(1'b0)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  rankings__m_axi
  (
    .clk(ap_clk),
    .rst(rankings__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_rankings_ARADDR),
    .m_axi_ARBURST(m_axi_rankings_ARBURST),
    .m_axi_ARCACHE(m_axi_rankings_ARCACHE),
    .m_axi_ARID(m_axi_rankings_ARID),
    .m_axi_ARLEN(m_axi_rankings_ARLEN),
    .m_axi_ARLOCK(m_axi_rankings_ARLOCK),
    .m_axi_ARPROT(m_axi_rankings_ARPROT),
    .m_axi_ARQOS(m_axi_rankings_ARQOS),
    .m_axi_ARREADY(m_axi_rankings_ARREADY),
    .m_axi_ARREGION(m_axi_rankings_ARREGION),
    .m_axi_ARSIZE(m_axi_rankings_ARSIZE),
    .m_axi_ARUSER(m_axi_rankings_ARUSER),
    .m_axi_ARVALID(m_axi_rankings_ARVALID),
    .m_axi_AWADDR(m_axi_rankings_AWADDR),
    .m_axi_AWBURST(m_axi_rankings_AWBURST),
    .m_axi_AWCACHE(m_axi_rankings_AWCACHE),
    .m_axi_AWID(m_axi_rankings_AWID),
    .m_axi_AWLEN(m_axi_rankings_AWLEN),
    .m_axi_AWLOCK(m_axi_rankings_AWLOCK),
    .m_axi_AWPROT(m_axi_rankings_AWPROT),
    .m_axi_AWQOS(m_axi_rankings_AWQOS),
    .m_axi_AWREADY(m_axi_rankings_AWREADY),
    .m_axi_AWREGION(m_axi_rankings_AWREGION),
    .m_axi_AWSIZE(m_axi_rankings_AWSIZE),
    .m_axi_AWUSER(m_axi_rankings_AWUSER),
    .m_axi_AWVALID(m_axi_rankings_AWVALID),
    .m_axi_BID(m_axi_rankings_BID),
    .m_axi_BREADY(m_axi_rankings_BREADY),
    .m_axi_BRESP(m_axi_rankings_BRESP),
    .m_axi_BUSER(m_axi_rankings_BUSER),
    .m_axi_BVALID(m_axi_rankings_BVALID),
    .m_axi_RDATA(m_axi_rankings_RDATA),
    .m_axi_RID(m_axi_rankings_RID),
    .m_axi_RLAST(m_axi_rankings_RLAST),
    .m_axi_RREADY(m_axi_rankings_RREADY),
    .m_axi_RRESP(m_axi_rankings_RRESP),
    .m_axi_RUSER(m_axi_rankings_RUSER),
    .m_axi_RVALID(m_axi_rankings_RVALID),
    .m_axi_WDATA(m_axi_rankings_WDATA),
    .m_axi_WID(m_axi_rankings_WID),
    .m_axi_WLAST(m_axi_rankings_WLAST),
    .m_axi_WREADY(m_axi_rankings_WREADY),
    .m_axi_WSTRB(m_axi_rankings_WSTRB),
    .m_axi_WUSER(m_axi_rankings_WUSER),
    .m_axi_WVALID(m_axi_rankings_WVALID),
    .read_addr_din(rankings__q2 + {rankings_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(rankings_read_addr__full_n),
    .read_addr_write(rankings_read_addr__write),
    .read_data_dout(rankings_read_data__dout),
    .read_data_empty_n(rankings_read_data__empty_n),
    .read_data_read(rankings_read_data__read),
    .write_addr_din(rankings__q2 + {rankings_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(rankings_write_addr__full_n),
    .write_addr_write(rankings_write_addr__write),
    .write_data_din(rankings_write_data__din),
    .write_data_full_n(rankings_write_data__full_n),
    .write_data_write(rankings_write_data__write)
  );


  async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .BurstLenWidth(3)
  )
  tmps__m_axi
  (
    .clk(ap_clk),
    .rst(tmps__rst__q2),
    .max_wait_time(2'd3),
    .max_burst_len(3'd7),
    .m_axi_ARADDR(m_axi_tmps_ARADDR),
    .m_axi_ARBURST(m_axi_tmps_ARBURST),
    .m_axi_ARCACHE(m_axi_tmps_ARCACHE),
    .m_axi_ARID(m_axi_tmps_ARID),
    .m_axi_ARLEN(m_axi_tmps_ARLEN),
    .m_axi_ARLOCK(m_axi_tmps_ARLOCK),
    .m_axi_ARPROT(m_axi_tmps_ARPROT),
    .m_axi_ARQOS(m_axi_tmps_ARQOS),
    .m_axi_ARREADY(m_axi_tmps_ARREADY),
    .m_axi_ARREGION(m_axi_tmps_ARREGION),
    .m_axi_ARSIZE(m_axi_tmps_ARSIZE),
    .m_axi_ARUSER(m_axi_tmps_ARUSER),
    .m_axi_ARVALID(m_axi_tmps_ARVALID),
    .m_axi_AWADDR(m_axi_tmps_AWADDR),
    .m_axi_AWBURST(m_axi_tmps_AWBURST),
    .m_axi_AWCACHE(m_axi_tmps_AWCACHE),
    .m_axi_AWID(m_axi_tmps_AWID),
    .m_axi_AWLEN(m_axi_tmps_AWLEN),
    .m_axi_AWLOCK(m_axi_tmps_AWLOCK),
    .m_axi_AWPROT(m_axi_tmps_AWPROT),
    .m_axi_AWQOS(m_axi_tmps_AWQOS),
    .m_axi_AWREADY(m_axi_tmps_AWREADY),
    .m_axi_AWREGION(m_axi_tmps_AWREGION),
    .m_axi_AWSIZE(m_axi_tmps_AWSIZE),
    .m_axi_AWUSER(m_axi_tmps_AWUSER),
    .m_axi_AWVALID(m_axi_tmps_AWVALID),
    .m_axi_BID(m_axi_tmps_BID),
    .m_axi_BREADY(m_axi_tmps_BREADY),
    .m_axi_BRESP(m_axi_tmps_BRESP),
    .m_axi_BUSER(m_axi_tmps_BUSER),
    .m_axi_BVALID(m_axi_tmps_BVALID),
    .m_axi_RDATA(m_axi_tmps_RDATA),
    .m_axi_RID(m_axi_tmps_RID),
    .m_axi_RLAST(m_axi_tmps_RLAST),
    .m_axi_RREADY(m_axi_tmps_RREADY),
    .m_axi_RRESP(m_axi_tmps_RRESP),
    .m_axi_RUSER(m_axi_tmps_RUSER),
    .m_axi_RVALID(m_axi_tmps_RVALID),
    .m_axi_WDATA(m_axi_tmps_WDATA),
    .m_axi_WID(m_axi_tmps_WID),
    .m_axi_WLAST(m_axi_tmps_WLAST),
    .m_axi_WREADY(m_axi_tmps_WREADY),
    .m_axi_WSTRB(m_axi_tmps_WSTRB),
    .m_axi_WUSER(m_axi_tmps_WUSER),
    .m_axi_WVALID(m_axi_tmps_WVALID),
    .read_addr_din(tmps__q2 + {tmps_read_addr__din[57:0], 6'd0}),
    .read_addr_full_n(tmps_read_addr__full_n),
    .read_addr_write(tmps_read_addr__write),
    .read_data_dout(tmps_read_data__dout),
    .read_data_empty_n(tmps_read_data__empty_n),
    .read_data_read(tmps_read_data__read),
    .write_addr_din(tmps__q2 + {tmps_write_addr__din[57:0], 6'd0}),
    .write_addr_full_n(tmps_write_addr__full_n),
    .write_addr_write(tmps_write_addr__write),
    .write_data_din(tmps_write_data__din),
    .write_data_full_n(tmps_write_data__full_n),
    .write_data_write(tmps_write_data__write)
  );


  always @(posedge ap_clk) begin
    ap_rst_n__q1 <= ap_rst_n__q0;
    ap_rst_n__q2 <= ap_rst_n__q1;
  end

  assign ap_rst_n__q0 = ap_rst_n;
  assign ap_rst_n_inv = (~ap_rst_n__q2);

  always @(posedge ap_clk) begin
    edge_req_0__rst__q1 <= edge_req_0__rst__q0;
    edge_req_0__rst__q2 <= edge_req_0__rst__q1;
  end

  assign edge_req_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_req_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             edge_req[0]\033[0m -> \033[90mEdgeMem_0               \033[0m %h", edge_req_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_req_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_0\033[0m -> \033[97medge_req[0]             \033[0m %h", edge_req_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_req_1__rst__q1 <= edge_req_1__rst__q0;
    edge_req_1__rst__q2 <= edge_req_1__rst__q1;
  end

  assign edge_req_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_req_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             edge_req[1]\033[0m -> \033[90mEdgeMem_1               \033[0m %h", edge_req_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_req_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_1\033[0m -> \033[97medge_req[1]             \033[0m %h", edge_req_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_req_2__rst__q1 <= edge_req_2__rst__q0;
    edge_req_2__rst__q2 <= edge_req_2__rst__q1;
  end

  assign edge_req_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_req_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             edge_req[2]\033[0m -> \033[90mEdgeMem_2               \033[0m %h", edge_req_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_req_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_2\033[0m -> \033[97medge_req[2]             \033[0m %h", edge_req_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_req_3__rst__q1 <= edge_req_3__rst__q0;
    edge_req_3__rst__q2 <= edge_req_3__rst__q1;
  end

  assign edge_req_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_req_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             edge_req[3]\033[0m -> \033[90mEdgeMem_3               \033[0m %h", edge_req_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_req_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_3\033[0m -> \033[97medge_req[3]             \033[0m %h", edge_req_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_req_4__rst__q1 <= edge_req_4__rst__q0;
    edge_req_4__rst__q2 <= edge_req_4__rst__q1;
  end

  assign edge_req_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_req_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             edge_req[4]\033[0m -> \033[90mEdgeMem_4               \033[0m %h", edge_req_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_req_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_4\033[0m -> \033[97medge_req[4]             \033[0m %h", edge_req_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_req_5__rst__q1 <= edge_req_5__rst__q0;
    edge_req_5__rst__q2 <= edge_req_5__rst__q1;
  end

  assign edge_req_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_req_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             edge_req[5]\033[0m -> \033[90mEdgeMem_5               \033[0m %h", edge_req_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_req_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_5\033[0m -> \033[97medge_req[5]             \033[0m %h", edge_req_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_req_6__rst__q1 <= edge_req_6__rst__q0;
    edge_req_6__rst__q2 <= edge_req_6__rst__q1;
  end

  assign edge_req_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_req_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             edge_req[6]\033[0m -> \033[90mEdgeMem_6               \033[0m %h", edge_req_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_req_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_6\033[0m -> \033[97medge_req[6]             \033[0m %h", edge_req_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_req_7__rst__q1 <= edge_req_7__rst__q0;
    edge_req_7__rst__q2 <= edge_req_7__rst__q1;
  end

  assign edge_req_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_req_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             edge_req[7]\033[0m -> \033[90mEdgeMem_7               \033[0m %h", edge_req_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_req_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_7\033[0m -> \033[97medge_req[7]             \033[0m %h", edge_req_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_resp_0__rst__q1 <= edge_resp_0__rst__q0;
    edge_resp_0__rst__q2 <= edge_resp_0__rst__q1;
  end

  assign edge_resp_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_resp_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            edge_resp[0]\033[0m -> \033[90mProcElem_0              \033[0m %h", edge_resp_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_resp_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               EdgeMem_0\033[0m -> \033[97medge_resp[0]            \033[0m %h", edge_resp_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_resp_1__rst__q1 <= edge_resp_1__rst__q0;
    edge_resp_1__rst__q2 <= edge_resp_1__rst__q1;
  end

  assign edge_resp_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_resp_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            edge_resp[1]\033[0m -> \033[90mProcElem_1              \033[0m %h", edge_resp_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_resp_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               EdgeMem_1\033[0m -> \033[97medge_resp[1]            \033[0m %h", edge_resp_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_resp_2__rst__q1 <= edge_resp_2__rst__q0;
    edge_resp_2__rst__q2 <= edge_resp_2__rst__q1;
  end

  assign edge_resp_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_resp_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            edge_resp[2]\033[0m -> \033[90mProcElem_2              \033[0m %h", edge_resp_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_resp_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               EdgeMem_2\033[0m -> \033[97medge_resp[2]            \033[0m %h", edge_resp_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_resp_3__rst__q1 <= edge_resp_3__rst__q0;
    edge_resp_3__rst__q2 <= edge_resp_3__rst__q1;
  end

  assign edge_resp_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_resp_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            edge_resp[3]\033[0m -> \033[90mProcElem_3              \033[0m %h", edge_resp_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_resp_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               EdgeMem_3\033[0m -> \033[97medge_resp[3]            \033[0m %h", edge_resp_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_resp_4__rst__q1 <= edge_resp_4__rst__q0;
    edge_resp_4__rst__q2 <= edge_resp_4__rst__q1;
  end

  assign edge_resp_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_resp_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            edge_resp[4]\033[0m -> \033[90mProcElem_4              \033[0m %h", edge_resp_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_resp_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               EdgeMem_4\033[0m -> \033[97medge_resp[4]            \033[0m %h", edge_resp_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_resp_5__rst__q1 <= edge_resp_5__rst__q0;
    edge_resp_5__rst__q2 <= edge_resp_5__rst__q1;
  end

  assign edge_resp_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_resp_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            edge_resp[5]\033[0m -> \033[90mProcElem_5              \033[0m %h", edge_resp_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_resp_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               EdgeMem_5\033[0m -> \033[97medge_resp[5]            \033[0m %h", edge_resp_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_resp_6__rst__q1 <= edge_resp_6__rst__q0;
    edge_resp_6__rst__q2 <= edge_resp_6__rst__q1;
  end

  assign edge_resp_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_resp_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            edge_resp[6]\033[0m -> \033[90mProcElem_6              \033[0m %h", edge_resp_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_resp_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               EdgeMem_6\033[0m -> \033[97medge_resp[6]            \033[0m %h", edge_resp_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    edge_resp_7__rst__q1 <= edge_resp_7__rst__q0;
    edge_resp_7__rst__q2 <= edge_resp_7__rst__q1;
  end

  assign edge_resp_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(edge_resp_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            edge_resp[7]\033[0m -> \033[90mProcElem_7              \033[0m %h", edge_resp_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(edge_resp_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               EdgeMem_7\033[0m -> \033[97medge_resp[7]            \033[0m %h", edge_resp_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    num_updates_0__rst__q1 <= num_updates_0__rst__q0;
    num_updates_0__rst__q2 <= num_updates_0__rst__q1;
  end

  assign num_updates_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(num_updates_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m          num_updates[0]\033[0m -> \033[90mControl_0               \033[0m %h", num_updates_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(num_updates_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_0\033[0m -> \033[97mnum_updates[0]          \033[0m %h", num_updates_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    num_updates_1__rst__q1 <= num_updates_1__rst__q0;
    num_updates_1__rst__q2 <= num_updates_1__rst__q1;
  end

  assign num_updates_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(num_updates_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m          num_updates[1]\033[0m -> \033[90mControl_0               \033[0m %h", num_updates_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(num_updates_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_1\033[0m -> \033[97mnum_updates[1]          \033[0m %h", num_updates_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    num_updates_2__rst__q1 <= num_updates_2__rst__q0;
    num_updates_2__rst__q2 <= num_updates_2__rst__q1;
  end

  assign num_updates_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(num_updates_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m          num_updates[2]\033[0m -> \033[90mControl_0               \033[0m %h", num_updates_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(num_updates_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_2\033[0m -> \033[97mnum_updates[2]          \033[0m %h", num_updates_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    num_updates_3__rst__q1 <= num_updates_3__rst__q0;
    num_updates_3__rst__q2 <= num_updates_3__rst__q1;
  end

  assign num_updates_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(num_updates_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m          num_updates[3]\033[0m -> \033[90mControl_0               \033[0m %h", num_updates_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(num_updates_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_3\033[0m -> \033[97mnum_updates[3]          \033[0m %h", num_updates_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    num_updates_4__rst__q1 <= num_updates_4__rst__q0;
    num_updates_4__rst__q2 <= num_updates_4__rst__q1;
  end

  assign num_updates_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(num_updates_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m          num_updates[4]\033[0m -> \033[90mControl_0               \033[0m %h", num_updates_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(num_updates_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_4\033[0m -> \033[97mnum_updates[4]          \033[0m %h", num_updates_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    num_updates_5__rst__q1 <= num_updates_5__rst__q0;
    num_updates_5__rst__q2 <= num_updates_5__rst__q1;
  end

  assign num_updates_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(num_updates_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m          num_updates[5]\033[0m -> \033[90mControl_0               \033[0m %h", num_updates_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(num_updates_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_5\033[0m -> \033[97mnum_updates[5]          \033[0m %h", num_updates_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    num_updates_6__rst__q1 <= num_updates_6__rst__q0;
    num_updates_6__rst__q2 <= num_updates_6__rst__q1;
  end

  assign num_updates_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(num_updates_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m          num_updates[6]\033[0m -> \033[90mControl_0               \033[0m %h", num_updates_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(num_updates_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_6\033[0m -> \033[97mnum_updates[6]          \033[0m %h", num_updates_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    num_updates_7__rst__q1 <= num_updates_7__rst__q0;
    num_updates_7__rst__q2 <= num_updates_7__rst__q1;
  end

  assign num_updates_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(num_updates_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m          num_updates[7]\033[0m -> \033[90mControl_0               \033[0m %h", num_updates_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(num_updates_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_7\033[0m -> \033[97mnum_updates[7]          \033[0m %h", num_updates_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    scatter_phase_vertex_req__rst__q1 <= scatter_phase_vertex_req__rst__q0;
    scatter_phase_vertex_req__rst__q2 <= scatter_phase_vertex_req__rst__q1;
  end

  assign scatter_phase_vertex_req__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(scatter_phase_vertex_req__read == 1'b1) begin
      $display("DEBUG: R: \033[97mscatter_phase_vertex_req\033[0m -> \033[90mVertexMem_0             \033[0m %h", scatter_phase_vertex_req__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(scatter_phase_vertex_req__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mscatter_phase_vertex_req\033[0m %h", scatter_phase_vertex_req__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_req_0__rst__q1 <= task_req_0__rst__q0;
    task_req_0__rst__q2 <= task_req_0__rst__q1;
  end

  assign task_req_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_req_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             task_req[0]\033[0m -> \033[90mProcElem_0              \033[0m %h", task_req_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_req_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mtask_req[0]             \033[0m %h", task_req_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_req_1__rst__q1 <= task_req_1__rst__q0;
    task_req_1__rst__q2 <= task_req_1__rst__q1;
  end

  assign task_req_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_req_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             task_req[1]\033[0m -> \033[90mProcElem_1              \033[0m %h", task_req_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_req_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mtask_req[1]             \033[0m %h", task_req_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_req_2__rst__q1 <= task_req_2__rst__q0;
    task_req_2__rst__q2 <= task_req_2__rst__q1;
  end

  assign task_req_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_req_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             task_req[2]\033[0m -> \033[90mProcElem_2              \033[0m %h", task_req_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_req_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mtask_req[2]             \033[0m %h", task_req_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_req_3__rst__q1 <= task_req_3__rst__q0;
    task_req_3__rst__q2 <= task_req_3__rst__q1;
  end

  assign task_req_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_req_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             task_req[3]\033[0m -> \033[90mProcElem_3              \033[0m %h", task_req_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_req_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mtask_req[3]             \033[0m %h", task_req_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_req_4__rst__q1 <= task_req_4__rst__q0;
    task_req_4__rst__q2 <= task_req_4__rst__q1;
  end

  assign task_req_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_req_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             task_req[4]\033[0m -> \033[90mProcElem_4              \033[0m %h", task_req_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_req_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mtask_req[4]             \033[0m %h", task_req_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_req_5__rst__q1 <= task_req_5__rst__q0;
    task_req_5__rst__q2 <= task_req_5__rst__q1;
  end

  assign task_req_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_req_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             task_req[5]\033[0m -> \033[90mProcElem_5              \033[0m %h", task_req_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_req_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mtask_req[5]             \033[0m %h", task_req_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_req_6__rst__q1 <= task_req_6__rst__q0;
    task_req_6__rst__q2 <= task_req_6__rst__q1;
  end

  assign task_req_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_req_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             task_req[6]\033[0m -> \033[90mProcElem_6              \033[0m %h", task_req_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_req_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mtask_req[6]             \033[0m %h", task_req_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_req_7__rst__q1 <= task_req_7__rst__q0;
    task_req_7__rst__q2 <= task_req_7__rst__q1;
  end

  assign task_req_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_req_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m             task_req[7]\033[0m -> \033[90mProcElem_7              \033[0m %h", task_req_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_req_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mtask_req[7]             \033[0m %h", task_req_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_resp_0__rst__q1 <= task_resp_0__rst__q0;
    task_resp_0__rst__q2 <= task_resp_0__rst__q1;
  end

  assign task_resp_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_resp_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            task_resp[0]\033[0m -> \033[90mControl_0               \033[0m %h", task_resp_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_resp_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_0\033[0m -> \033[97mtask_resp[0]            \033[0m %h", task_resp_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_resp_1__rst__q1 <= task_resp_1__rst__q0;
    task_resp_1__rst__q2 <= task_resp_1__rst__q1;
  end

  assign task_resp_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_resp_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            task_resp[1]\033[0m -> \033[90mControl_0               \033[0m %h", task_resp_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_resp_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_1\033[0m -> \033[97mtask_resp[1]            \033[0m %h", task_resp_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_resp_2__rst__q1 <= task_resp_2__rst__q0;
    task_resp_2__rst__q2 <= task_resp_2__rst__q1;
  end

  assign task_resp_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_resp_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            task_resp[2]\033[0m -> \033[90mControl_0               \033[0m %h", task_resp_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_resp_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_2\033[0m -> \033[97mtask_resp[2]            \033[0m %h", task_resp_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_resp_3__rst__q1 <= task_resp_3__rst__q0;
    task_resp_3__rst__q2 <= task_resp_3__rst__q1;
  end

  assign task_resp_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_resp_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            task_resp[3]\033[0m -> \033[90mControl_0               \033[0m %h", task_resp_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_resp_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_3\033[0m -> \033[97mtask_resp[3]            \033[0m %h", task_resp_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_resp_4__rst__q1 <= task_resp_4__rst__q0;
    task_resp_4__rst__q2 <= task_resp_4__rst__q1;
  end

  assign task_resp_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_resp_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            task_resp[4]\033[0m -> \033[90mControl_0               \033[0m %h", task_resp_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_resp_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_4\033[0m -> \033[97mtask_resp[4]            \033[0m %h", task_resp_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_resp_5__rst__q1 <= task_resp_5__rst__q0;
    task_resp_5__rst__q2 <= task_resp_5__rst__q1;
  end

  assign task_resp_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_resp_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            task_resp[5]\033[0m -> \033[90mControl_0               \033[0m %h", task_resp_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_resp_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_5\033[0m -> \033[97mtask_resp[5]            \033[0m %h", task_resp_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_resp_6__rst__q1 <= task_resp_6__rst__q0;
    task_resp_6__rst__q2 <= task_resp_6__rst__q1;
  end

  assign task_resp_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_resp_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            task_resp[6]\033[0m -> \033[90mControl_0               \033[0m %h", task_resp_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_resp_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_6\033[0m -> \033[97mtask_resp[6]            \033[0m %h", task_resp_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    task_resp_7__rst__q1 <= task_resp_7__rst__q0;
    task_resp_7__rst__q2 <= task_resp_7__rst__q1;
  end

  assign task_resp_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(task_resp_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m            task_resp[7]\033[0m -> \033[90mControl_0               \033[0m %h", task_resp_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(task_resp_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_7\033[0m -> \033[97mtask_resp[7]            \033[0m %h", task_resp_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_config_0__rst__q1 <= update_config_0__rst__q0;
    update_config_0__rst__q2 <= update_config_0__rst__q1;
  end

  assign update_config_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_config_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        update_config[0]\033[0m -> \033[90mUpdateHandler_0         \033[0m %h", update_config_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_config_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_config[0]        \033[0m %h", update_config_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_config_1__rst__q1 <= update_config_1__rst__q0;
    update_config_1__rst__q2 <= update_config_1__rst__q1;
  end

  assign update_config_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_config_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        update_config[1]\033[0m -> \033[90mUpdateHandler_1         \033[0m %h", update_config_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_config_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_config[1]        \033[0m %h", update_config_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_config_2__rst__q1 <= update_config_2__rst__q0;
    update_config_2__rst__q2 <= update_config_2__rst__q1;
  end

  assign update_config_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_config_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        update_config[2]\033[0m -> \033[90mUpdateHandler_2         \033[0m %h", update_config_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_config_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_config[2]        \033[0m %h", update_config_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_config_3__rst__q1 <= update_config_3__rst__q0;
    update_config_3__rst__q2 <= update_config_3__rst__q1;
  end

  assign update_config_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_config_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        update_config[3]\033[0m -> \033[90mUpdateHandler_3         \033[0m %h", update_config_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_config_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_config[3]        \033[0m %h", update_config_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_config_4__rst__q1 <= update_config_4__rst__q0;
    update_config_4__rst__q2 <= update_config_4__rst__q1;
  end

  assign update_config_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_config_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        update_config[4]\033[0m -> \033[90mUpdateHandler_4         \033[0m %h", update_config_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_config_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_config[4]        \033[0m %h", update_config_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_config_5__rst__q1 <= update_config_5__rst__q0;
    update_config_5__rst__q2 <= update_config_5__rst__q1;
  end

  assign update_config_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_config_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        update_config[5]\033[0m -> \033[90mUpdateHandler_5         \033[0m %h", update_config_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_config_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_config[5]        \033[0m %h", update_config_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_config_6__rst__q1 <= update_config_6__rst__q0;
    update_config_6__rst__q2 <= update_config_6__rst__q1;
  end

  assign update_config_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_config_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        update_config[6]\033[0m -> \033[90mUpdateHandler_6         \033[0m %h", update_config_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_config_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_config[6]        \033[0m %h", update_config_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_config_7__rst__q1 <= update_config_7__rst__q0;
    update_config_7__rst__q2 <= update_config_7__rst__q1;
  end

  assign update_config_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_config_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        update_config[7]\033[0m -> \033[90mUpdateHandler_7         \033[0m %h", update_config_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_config_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_config[7]        \033[0m %h", update_config_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_mm2pe_0__rst__q1 <= update_mm2pe_0__rst__q0;
    update_mm2pe_0__rst__q2 <= update_mm2pe_0__rst__q1;
  end

  assign update_mm2pe_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_mm2pe_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_mm2pe[0]\033[0m -> \033[90mProcElem_0              \033[0m %h", update_mm2pe_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_mm2pe_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_0\033[0m -> \033[97mupdate_mm2pe[0]         \033[0m %h", update_mm2pe_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_mm2pe_1__rst__q1 <= update_mm2pe_1__rst__q0;
    update_mm2pe_1__rst__q2 <= update_mm2pe_1__rst__q1;
  end

  assign update_mm2pe_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_mm2pe_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_mm2pe[1]\033[0m -> \033[90mProcElem_1              \033[0m %h", update_mm2pe_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_mm2pe_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_1\033[0m -> \033[97mupdate_mm2pe[1]         \033[0m %h", update_mm2pe_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_mm2pe_2__rst__q1 <= update_mm2pe_2__rst__q0;
    update_mm2pe_2__rst__q2 <= update_mm2pe_2__rst__q1;
  end

  assign update_mm2pe_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_mm2pe_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_mm2pe[2]\033[0m -> \033[90mProcElem_2              \033[0m %h", update_mm2pe_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_mm2pe_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_2\033[0m -> \033[97mupdate_mm2pe[2]         \033[0m %h", update_mm2pe_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_mm2pe_3__rst__q1 <= update_mm2pe_3__rst__q0;
    update_mm2pe_3__rst__q2 <= update_mm2pe_3__rst__q1;
  end

  assign update_mm2pe_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_mm2pe_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_mm2pe[3]\033[0m -> \033[90mProcElem_3              \033[0m %h", update_mm2pe_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_mm2pe_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_3\033[0m -> \033[97mupdate_mm2pe[3]         \033[0m %h", update_mm2pe_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_mm2pe_4__rst__q1 <= update_mm2pe_4__rst__q0;
    update_mm2pe_4__rst__q2 <= update_mm2pe_4__rst__q1;
  end

  assign update_mm2pe_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_mm2pe_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_mm2pe[4]\033[0m -> \033[90mProcElem_4              \033[0m %h", update_mm2pe_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_mm2pe_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_4\033[0m -> \033[97mupdate_mm2pe[4]         \033[0m %h", update_mm2pe_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_mm2pe_5__rst__q1 <= update_mm2pe_5__rst__q0;
    update_mm2pe_5__rst__q2 <= update_mm2pe_5__rst__q1;
  end

  assign update_mm2pe_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_mm2pe_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_mm2pe[5]\033[0m -> \033[90mProcElem_5              \033[0m %h", update_mm2pe_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_mm2pe_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_5\033[0m -> \033[97mupdate_mm2pe[5]         \033[0m %h", update_mm2pe_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_mm2pe_6__rst__q1 <= update_mm2pe_6__rst__q0;
    update_mm2pe_6__rst__q2 <= update_mm2pe_6__rst__q1;
  end

  assign update_mm2pe_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_mm2pe_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_mm2pe[6]\033[0m -> \033[90mProcElem_6              \033[0m %h", update_mm2pe_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_mm2pe_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_6\033[0m -> \033[97mupdate_mm2pe[6]         \033[0m %h", update_mm2pe_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_mm2pe_7__rst__q1 <= update_mm2pe_7__rst__q0;
    update_mm2pe_7__rst__q2 <= update_mm2pe_7__rst__q1;
  end

  assign update_mm2pe_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_mm2pe_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_mm2pe[7]\033[0m -> \033[90mProcElem_7              \033[0m %h", update_mm2pe_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_mm2pe_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_7\033[0m -> \033[97mupdate_mm2pe[7]         \033[0m %h", update_mm2pe_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_pe2mm_0__rst__q1 <= update_pe2mm_0__rst__q0;
    update_pe2mm_0__rst__q2 <= update_pe2mm_0__rst__q1;
  end

  assign update_pe2mm_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_pe2mm_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_pe2mm[0]\033[0m -> \033[90mUpdateHandler_0         \033[0m %h", update_pe2mm_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_pe2mm_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_0\033[0m -> \033[97mupdate_pe2mm[0]         \033[0m %h", update_pe2mm_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_pe2mm_1__rst__q1 <= update_pe2mm_1__rst__q0;
    update_pe2mm_1__rst__q2 <= update_pe2mm_1__rst__q1;
  end

  assign update_pe2mm_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_pe2mm_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_pe2mm[1]\033[0m -> \033[90mUpdateHandler_1         \033[0m %h", update_pe2mm_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_pe2mm_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_1\033[0m -> \033[97mupdate_pe2mm[1]         \033[0m %h", update_pe2mm_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_pe2mm_2__rst__q1 <= update_pe2mm_2__rst__q0;
    update_pe2mm_2__rst__q2 <= update_pe2mm_2__rst__q1;
  end

  assign update_pe2mm_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_pe2mm_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_pe2mm[2]\033[0m -> \033[90mUpdateHandler_2         \033[0m %h", update_pe2mm_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_pe2mm_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_2\033[0m -> \033[97mupdate_pe2mm[2]         \033[0m %h", update_pe2mm_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_pe2mm_3__rst__q1 <= update_pe2mm_3__rst__q0;
    update_pe2mm_3__rst__q2 <= update_pe2mm_3__rst__q1;
  end

  assign update_pe2mm_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_pe2mm_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_pe2mm[3]\033[0m -> \033[90mUpdateHandler_3         \033[0m %h", update_pe2mm_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_pe2mm_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_3\033[0m -> \033[97mupdate_pe2mm[3]         \033[0m %h", update_pe2mm_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_pe2mm_4__rst__q1 <= update_pe2mm_4__rst__q0;
    update_pe2mm_4__rst__q2 <= update_pe2mm_4__rst__q1;
  end

  assign update_pe2mm_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_pe2mm_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_pe2mm[4]\033[0m -> \033[90mUpdateHandler_4         \033[0m %h", update_pe2mm_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_pe2mm_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_4\033[0m -> \033[97mupdate_pe2mm[4]         \033[0m %h", update_pe2mm_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_pe2mm_5__rst__q1 <= update_pe2mm_5__rst__q0;
    update_pe2mm_5__rst__q2 <= update_pe2mm_5__rst__q1;
  end

  assign update_pe2mm_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_pe2mm_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_pe2mm[5]\033[0m -> \033[90mUpdateHandler_5         \033[0m %h", update_pe2mm_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_pe2mm_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_5\033[0m -> \033[97mupdate_pe2mm[5]         \033[0m %h", update_pe2mm_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_pe2mm_6__rst__q1 <= update_pe2mm_6__rst__q0;
    update_pe2mm_6__rst__q2 <= update_pe2mm_6__rst__q1;
  end

  assign update_pe2mm_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_pe2mm_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_pe2mm[6]\033[0m -> \033[90mUpdateHandler_6         \033[0m %h", update_pe2mm_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_pe2mm_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_6\033[0m -> \033[97mupdate_pe2mm[6]         \033[0m %h", update_pe2mm_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_pe2mm_7__rst__q1 <= update_pe2mm_7__rst__q0;
    update_pe2mm_7__rst__q2 <= update_pe2mm_7__rst__q1;
  end

  assign update_pe2mm_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_pe2mm_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_pe2mm[7]\033[0m -> \033[90mUpdateHandler_7         \033[0m %h", update_pe2mm_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_pe2mm_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_7\033[0m -> \033[97mupdate_pe2mm[7]         \033[0m %h", update_pe2mm_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_phase_0__rst__q1 <= update_phase_0__rst__q0;
    update_phase_0__rst__q2 <= update_phase_0__rst__q1;
  end

  assign update_phase_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_phase_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_phase[0]\033[0m -> \033[90mUpdateHandler_0         \033[0m %h", update_phase_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_phase_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_phase[0]         \033[0m %h", update_phase_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_phase_1__rst__q1 <= update_phase_1__rst__q0;
    update_phase_1__rst__q2 <= update_phase_1__rst__q1;
  end

  assign update_phase_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_phase_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_phase[1]\033[0m -> \033[90mUpdateHandler_1         \033[0m %h", update_phase_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_phase_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_phase[1]         \033[0m %h", update_phase_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_phase_2__rst__q1 <= update_phase_2__rst__q0;
    update_phase_2__rst__q2 <= update_phase_2__rst__q1;
  end

  assign update_phase_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_phase_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_phase[2]\033[0m -> \033[90mUpdateHandler_2         \033[0m %h", update_phase_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_phase_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_phase[2]         \033[0m %h", update_phase_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_phase_3__rst__q1 <= update_phase_3__rst__q0;
    update_phase_3__rst__q2 <= update_phase_3__rst__q1;
  end

  assign update_phase_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_phase_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_phase[3]\033[0m -> \033[90mUpdateHandler_3         \033[0m %h", update_phase_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_phase_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_phase[3]         \033[0m %h", update_phase_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_phase_4__rst__q1 <= update_phase_4__rst__q0;
    update_phase_4__rst__q2 <= update_phase_4__rst__q1;
  end

  assign update_phase_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_phase_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_phase[4]\033[0m -> \033[90mUpdateHandler_4         \033[0m %h", update_phase_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_phase_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_phase[4]         \033[0m %h", update_phase_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_phase_5__rst__q1 <= update_phase_5__rst__q0;
    update_phase_5__rst__q2 <= update_phase_5__rst__q1;
  end

  assign update_phase_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_phase_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_phase[5]\033[0m -> \033[90mUpdateHandler_5         \033[0m %h", update_phase_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_phase_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_phase[5]         \033[0m %h", update_phase_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_phase_6__rst__q1 <= update_phase_6__rst__q0;
    update_phase_6__rst__q2 <= update_phase_6__rst__q1;
  end

  assign update_phase_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_phase_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_phase[6]\033[0m -> \033[90mUpdateHandler_6         \033[0m %h", update_phase_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_phase_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_phase[6]         \033[0m %h", update_phase_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_phase_7__rst__q1 <= update_phase_7__rst__q0;
    update_phase_7__rst__q2 <= update_phase_7__rst__q1;
  end

  assign update_phase_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_phase_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m         update_phase[7]\033[0m -> \033[90mUpdateHandler_7         \033[0m %h", update_phase_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_phase_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m               Control_0\033[0m -> \033[97mupdate_phase[7]         \033[0m %h", update_phase_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_addr_0__rst__q1 <= update_read_addr_0__rst__q0;
    update_read_addr_0__rst__q2 <= update_read_addr_0__rst__q1;
  end

  assign update_read_addr_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_addr_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_addr[0]\033[0m -> \033[90mUpdateMem_0             \033[0m %h", update_read_addr_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_addr_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_0\033[0m -> \033[97mupdate_read_addr[0]     \033[0m %h", update_read_addr_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_addr_1__rst__q1 <= update_read_addr_1__rst__q0;
    update_read_addr_1__rst__q2 <= update_read_addr_1__rst__q1;
  end

  assign update_read_addr_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_addr_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_addr[1]\033[0m -> \033[90mUpdateMem_1             \033[0m %h", update_read_addr_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_addr_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_1\033[0m -> \033[97mupdate_read_addr[1]     \033[0m %h", update_read_addr_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_addr_2__rst__q1 <= update_read_addr_2__rst__q0;
    update_read_addr_2__rst__q2 <= update_read_addr_2__rst__q1;
  end

  assign update_read_addr_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_addr_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_addr[2]\033[0m -> \033[90mUpdateMem_2             \033[0m %h", update_read_addr_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_addr_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_2\033[0m -> \033[97mupdate_read_addr[2]     \033[0m %h", update_read_addr_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_addr_3__rst__q1 <= update_read_addr_3__rst__q0;
    update_read_addr_3__rst__q2 <= update_read_addr_3__rst__q1;
  end

  assign update_read_addr_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_addr_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_addr[3]\033[0m -> \033[90mUpdateMem_3             \033[0m %h", update_read_addr_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_addr_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_3\033[0m -> \033[97mupdate_read_addr[3]     \033[0m %h", update_read_addr_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_addr_4__rst__q1 <= update_read_addr_4__rst__q0;
    update_read_addr_4__rst__q2 <= update_read_addr_4__rst__q1;
  end

  assign update_read_addr_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_addr_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_addr[4]\033[0m -> \033[90mUpdateMem_4             \033[0m %h", update_read_addr_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_addr_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_4\033[0m -> \033[97mupdate_read_addr[4]     \033[0m %h", update_read_addr_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_addr_5__rst__q1 <= update_read_addr_5__rst__q0;
    update_read_addr_5__rst__q2 <= update_read_addr_5__rst__q1;
  end

  assign update_read_addr_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_addr_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_addr[5]\033[0m -> \033[90mUpdateMem_5             \033[0m %h", update_read_addr_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_addr_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_5\033[0m -> \033[97mupdate_read_addr[5]     \033[0m %h", update_read_addr_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_addr_6__rst__q1 <= update_read_addr_6__rst__q0;
    update_read_addr_6__rst__q2 <= update_read_addr_6__rst__q1;
  end

  assign update_read_addr_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_addr_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_addr[6]\033[0m -> \033[90mUpdateMem_6             \033[0m %h", update_read_addr_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_addr_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_6\033[0m -> \033[97mupdate_read_addr[6]     \033[0m %h", update_read_addr_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_addr_7__rst__q1 <= update_read_addr_7__rst__q0;
    update_read_addr_7__rst__q2 <= update_read_addr_7__rst__q1;
  end

  assign update_read_addr_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_addr_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_addr[7]\033[0m -> \033[90mUpdateMem_7             \033[0m %h", update_read_addr_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_addr_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_7\033[0m -> \033[97mupdate_read_addr[7]     \033[0m %h", update_read_addr_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_data_0__rst__q1 <= update_read_data_0__rst__q0;
    update_read_data_0__rst__q2 <= update_read_data_0__rst__q1;
  end

  assign update_read_data_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_data_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_data[0]\033[0m -> \033[90mUpdateHandler_0         \033[0m %h", update_read_data_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_data_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             UpdateMem_0\033[0m -> \033[97mupdate_read_data[0]     \033[0m %h", update_read_data_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_data_1__rst__q1 <= update_read_data_1__rst__q0;
    update_read_data_1__rst__q2 <= update_read_data_1__rst__q1;
  end

  assign update_read_data_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_data_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_data[1]\033[0m -> \033[90mUpdateHandler_1         \033[0m %h", update_read_data_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_data_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             UpdateMem_1\033[0m -> \033[97mupdate_read_data[1]     \033[0m %h", update_read_data_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_data_2__rst__q1 <= update_read_data_2__rst__q0;
    update_read_data_2__rst__q2 <= update_read_data_2__rst__q1;
  end

  assign update_read_data_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_data_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_data[2]\033[0m -> \033[90mUpdateHandler_2         \033[0m %h", update_read_data_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_data_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             UpdateMem_2\033[0m -> \033[97mupdate_read_data[2]     \033[0m %h", update_read_data_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_data_3__rst__q1 <= update_read_data_3__rst__q0;
    update_read_data_3__rst__q2 <= update_read_data_3__rst__q1;
  end

  assign update_read_data_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_data_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_data[3]\033[0m -> \033[90mUpdateHandler_3         \033[0m %h", update_read_data_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_data_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             UpdateMem_3\033[0m -> \033[97mupdate_read_data[3]     \033[0m %h", update_read_data_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_data_4__rst__q1 <= update_read_data_4__rst__q0;
    update_read_data_4__rst__q2 <= update_read_data_4__rst__q1;
  end

  assign update_read_data_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_data_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_data[4]\033[0m -> \033[90mUpdateHandler_4         \033[0m %h", update_read_data_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_data_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             UpdateMem_4\033[0m -> \033[97mupdate_read_data[4]     \033[0m %h", update_read_data_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_data_5__rst__q1 <= update_read_data_5__rst__q0;
    update_read_data_5__rst__q2 <= update_read_data_5__rst__q1;
  end

  assign update_read_data_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_data_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_data[5]\033[0m -> \033[90mUpdateHandler_5         \033[0m %h", update_read_data_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_data_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             UpdateMem_5\033[0m -> \033[97mupdate_read_data[5]     \033[0m %h", update_read_data_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_data_6__rst__q1 <= update_read_data_6__rst__q0;
    update_read_data_6__rst__q2 <= update_read_data_6__rst__q1;
  end

  assign update_read_data_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_data_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_data[6]\033[0m -> \033[90mUpdateHandler_6         \033[0m %h", update_read_data_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_data_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             UpdateMem_6\033[0m -> \033[97mupdate_read_data[6]     \033[0m %h", update_read_data_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_read_data_7__rst__q1 <= update_read_data_7__rst__q0;
    update_read_data_7__rst__q2 <= update_read_data_7__rst__q1;
  end

  assign update_read_data_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_read_data_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m     update_read_data[7]\033[0m -> \033[90mUpdateHandler_7         \033[0m %h", update_read_data_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_read_data_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             UpdateMem_7\033[0m -> \033[97mupdate_read_data[7]     \033[0m %h", update_read_data_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_req_0__rst__q1 <= update_req_0__rst__q0;
    update_req_0__rst__q2 <= update_req_0__rst__q1;
  end

  assign update_req_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_req_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m           update_req[0]\033[0m -> \033[90mUpdateHandler_0         \033[0m %h", update_req_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_req_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_0\033[0m -> \033[97mupdate_req[0]           \033[0m %h", update_req_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_req_1__rst__q1 <= update_req_1__rst__q0;
    update_req_1__rst__q2 <= update_req_1__rst__q1;
  end

  assign update_req_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_req_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m           update_req[1]\033[0m -> \033[90mUpdateHandler_1         \033[0m %h", update_req_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_req_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_1\033[0m -> \033[97mupdate_req[1]           \033[0m %h", update_req_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_req_2__rst__q1 <= update_req_2__rst__q0;
    update_req_2__rst__q2 <= update_req_2__rst__q1;
  end

  assign update_req_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_req_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m           update_req[2]\033[0m -> \033[90mUpdateHandler_2         \033[0m %h", update_req_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_req_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_2\033[0m -> \033[97mupdate_req[2]           \033[0m %h", update_req_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_req_3__rst__q1 <= update_req_3__rst__q0;
    update_req_3__rst__q2 <= update_req_3__rst__q1;
  end

  assign update_req_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_req_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m           update_req[3]\033[0m -> \033[90mUpdateHandler_3         \033[0m %h", update_req_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_req_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_3\033[0m -> \033[97mupdate_req[3]           \033[0m %h", update_req_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_req_4__rst__q1 <= update_req_4__rst__q0;
    update_req_4__rst__q2 <= update_req_4__rst__q1;
  end

  assign update_req_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_req_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m           update_req[4]\033[0m -> \033[90mUpdateHandler_4         \033[0m %h", update_req_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_req_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_4\033[0m -> \033[97mupdate_req[4]           \033[0m %h", update_req_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_req_5__rst__q1 <= update_req_5__rst__q0;
    update_req_5__rst__q2 <= update_req_5__rst__q1;
  end

  assign update_req_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_req_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m           update_req[5]\033[0m -> \033[90mUpdateHandler_5         \033[0m %h", update_req_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_req_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_5\033[0m -> \033[97mupdate_req[5]           \033[0m %h", update_req_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_req_6__rst__q1 <= update_req_6__rst__q0;
    update_req_6__rst__q2 <= update_req_6__rst__q1;
  end

  assign update_req_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_req_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m           update_req[6]\033[0m -> \033[90mUpdateHandler_6         \033[0m %h", update_req_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_req_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_6\033[0m -> \033[97mupdate_req[6]           \033[0m %h", update_req_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_req_7__rst__q1 <= update_req_7__rst__q0;
    update_req_7__rst__q2 <= update_req_7__rst__q1;
  end

  assign update_req_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_req_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m           update_req[7]\033[0m -> \033[90mUpdateHandler_7         \033[0m %h", update_req_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_req_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_7\033[0m -> \033[97mupdate_req[7]           \033[0m %h", update_req_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_addr_0__rst__q1 <= update_write_addr_0__rst__q0;
    update_write_addr_0__rst__q2 <= update_write_addr_0__rst__q1;
  end

  assign update_write_addr_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_addr_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_addr[0]\033[0m -> \033[90mUpdateMem_0             \033[0m %h", update_write_addr_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_addr_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_0\033[0m -> \033[97mupdate_write_addr[0]    \033[0m %h", update_write_addr_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_addr_1__rst__q1 <= update_write_addr_1__rst__q0;
    update_write_addr_1__rst__q2 <= update_write_addr_1__rst__q1;
  end

  assign update_write_addr_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_addr_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_addr[1]\033[0m -> \033[90mUpdateMem_1             \033[0m %h", update_write_addr_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_addr_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_1\033[0m -> \033[97mupdate_write_addr[1]    \033[0m %h", update_write_addr_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_addr_2__rst__q1 <= update_write_addr_2__rst__q0;
    update_write_addr_2__rst__q2 <= update_write_addr_2__rst__q1;
  end

  assign update_write_addr_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_addr_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_addr[2]\033[0m -> \033[90mUpdateMem_2             \033[0m %h", update_write_addr_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_addr_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_2\033[0m -> \033[97mupdate_write_addr[2]    \033[0m %h", update_write_addr_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_addr_3__rst__q1 <= update_write_addr_3__rst__q0;
    update_write_addr_3__rst__q2 <= update_write_addr_3__rst__q1;
  end

  assign update_write_addr_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_addr_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_addr[3]\033[0m -> \033[90mUpdateMem_3             \033[0m %h", update_write_addr_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_addr_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_3\033[0m -> \033[97mupdate_write_addr[3]    \033[0m %h", update_write_addr_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_addr_4__rst__q1 <= update_write_addr_4__rst__q0;
    update_write_addr_4__rst__q2 <= update_write_addr_4__rst__q1;
  end

  assign update_write_addr_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_addr_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_addr[4]\033[0m -> \033[90mUpdateMem_4             \033[0m %h", update_write_addr_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_addr_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_4\033[0m -> \033[97mupdate_write_addr[4]    \033[0m %h", update_write_addr_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_addr_5__rst__q1 <= update_write_addr_5__rst__q0;
    update_write_addr_5__rst__q2 <= update_write_addr_5__rst__q1;
  end

  assign update_write_addr_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_addr_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_addr[5]\033[0m -> \033[90mUpdateMem_5             \033[0m %h", update_write_addr_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_addr_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_5\033[0m -> \033[97mupdate_write_addr[5]    \033[0m %h", update_write_addr_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_addr_6__rst__q1 <= update_write_addr_6__rst__q0;
    update_write_addr_6__rst__q2 <= update_write_addr_6__rst__q1;
  end

  assign update_write_addr_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_addr_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_addr[6]\033[0m -> \033[90mUpdateMem_6             \033[0m %h", update_write_addr_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_addr_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_6\033[0m -> \033[97mupdate_write_addr[6]    \033[0m %h", update_write_addr_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_addr_7__rst__q1 <= update_write_addr_7__rst__q0;
    update_write_addr_7__rst__q2 <= update_write_addr_7__rst__q1;
  end

  assign update_write_addr_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_addr_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_addr[7]\033[0m -> \033[90mUpdateMem_7             \033[0m %h", update_write_addr_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_addr_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_7\033[0m -> \033[97mupdate_write_addr[7]    \033[0m %h", update_write_addr_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_data_0__rst__q1 <= update_write_data_0__rst__q0;
    update_write_data_0__rst__q2 <= update_write_data_0__rst__q1;
  end

  assign update_write_data_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_data_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_data[0]\033[0m -> \033[90mUpdateMem_0             \033[0m %h", update_write_data_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_data_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_0\033[0m -> \033[97mupdate_write_data[0]    \033[0m %h", update_write_data_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_data_1__rst__q1 <= update_write_data_1__rst__q0;
    update_write_data_1__rst__q2 <= update_write_data_1__rst__q1;
  end

  assign update_write_data_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_data_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_data[1]\033[0m -> \033[90mUpdateMem_1             \033[0m %h", update_write_data_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_data_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_1\033[0m -> \033[97mupdate_write_data[1]    \033[0m %h", update_write_data_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_data_2__rst__q1 <= update_write_data_2__rst__q0;
    update_write_data_2__rst__q2 <= update_write_data_2__rst__q1;
  end

  assign update_write_data_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_data_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_data[2]\033[0m -> \033[90mUpdateMem_2             \033[0m %h", update_write_data_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_data_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_2\033[0m -> \033[97mupdate_write_data[2]    \033[0m %h", update_write_data_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_data_3__rst__q1 <= update_write_data_3__rst__q0;
    update_write_data_3__rst__q2 <= update_write_data_3__rst__q1;
  end

  assign update_write_data_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_data_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_data[3]\033[0m -> \033[90mUpdateMem_3             \033[0m %h", update_write_data_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_data_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_3\033[0m -> \033[97mupdate_write_data[3]    \033[0m %h", update_write_data_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_data_4__rst__q1 <= update_write_data_4__rst__q0;
    update_write_data_4__rst__q2 <= update_write_data_4__rst__q1;
  end

  assign update_write_data_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_data_4__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_data[4]\033[0m -> \033[90mUpdateMem_4             \033[0m %h", update_write_data_4__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_data_4__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_4\033[0m -> \033[97mupdate_write_data[4]    \033[0m %h", update_write_data_4__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_data_5__rst__q1 <= update_write_data_5__rst__q0;
    update_write_data_5__rst__q2 <= update_write_data_5__rst__q1;
  end

  assign update_write_data_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_data_5__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_data[5]\033[0m -> \033[90mUpdateMem_5             \033[0m %h", update_write_data_5__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_data_5__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_5\033[0m -> \033[97mupdate_write_data[5]    \033[0m %h", update_write_data_5__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_data_6__rst__q1 <= update_write_data_6__rst__q0;
    update_write_data_6__rst__q2 <= update_write_data_6__rst__q1;
  end

  assign update_write_data_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_data_6__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_data[6]\033[0m -> \033[90mUpdateMem_6             \033[0m %h", update_write_data_6__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_data_6__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_6\033[0m -> \033[97mupdate_write_data[6]    \033[0m %h", update_write_data_6__din);
    end 
  end


  always @(posedge ap_clk) begin
    update_write_data_7__rst__q1 <= update_write_data_7__rst__q0;
    update_write_data_7__rst__q2 <= update_write_data_7__rst__q1;
  end

  assign update_write_data_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(update_write_data_7__read == 1'b1) begin
      $display("DEBUG: R: \033[97m    update_write_data[7]\033[0m -> \033[90mUpdateMem_7             \033[0m %h", update_write_data_7__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(update_write_data_7__write == 1'b1) begin
      $display("DEBUG: W: \033[90m         UpdateHandler_7\033[0m -> \033[97mupdate_write_data[7]    \033[0m %h", update_write_data_7__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r0_0__rst__q1 <= vertex_mm2pe_r0_0__rst__q0;
    vertex_mm2pe_r0_0__rst__q2 <= vertex_mm2pe_r0_0__rst__q1;
  end

  assign vertex_mm2pe_r0_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r0_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r0[0]\033[0m -> \033[90mProcElem_0              \033[0m %h", vertex_mm2pe_r0_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r0_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             VertexMem_0\033[0m -> \033[97mvertex_mm2pe_r0[0]      \033[0m %h", vertex_mm2pe_r0_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r0_1__rst__q1 <= vertex_mm2pe_r0_1__rst__q0;
    vertex_mm2pe_r0_1__rst__q2 <= vertex_mm2pe_r0_1__rst__q1;
  end

  assign vertex_mm2pe_r0_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r0_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r0[1]\033[0m -> \033[90mVertexRouterR1_0        \033[0m %h", vertex_mm2pe_r0_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r0_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m             VertexMem_0\033[0m -> \033[97mvertex_mm2pe_r0[1]      \033[0m %h", vertex_mm2pe_r0_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r1_0__rst__q1 <= vertex_mm2pe_r1_0__rst__q0;
    vertex_mm2pe_r1_0__rst__q2 <= vertex_mm2pe_r1_0__rst__q1;
  end

  assign vertex_mm2pe_r1_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r1_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r1[0]\033[0m -> \033[90mProcElem_1              \033[0m %h", vertex_mm2pe_r1_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r1_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR1_0\033[0m -> \033[97mvertex_mm2pe_r1[0]      \033[0m %h", vertex_mm2pe_r1_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r1_1__rst__q1 <= vertex_mm2pe_r1_1__rst__q0;
    vertex_mm2pe_r1_1__rst__q2 <= vertex_mm2pe_r1_1__rst__q1;
  end

  assign vertex_mm2pe_r1_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r1_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r1[1]\033[0m -> \033[90mProcElem_2              \033[0m %h", vertex_mm2pe_r1_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r1_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR1_0\033[0m -> \033[97mvertex_mm2pe_r1[1]      \033[0m %h", vertex_mm2pe_r1_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r1_2__rst__q1 <= vertex_mm2pe_r1_2__rst__q0;
    vertex_mm2pe_r1_2__rst__q2 <= vertex_mm2pe_r1_2__rst__q1;
  end

  assign vertex_mm2pe_r1_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r1_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r1[2]\033[0m -> \033[90mProcElem_3              \033[0m %h", vertex_mm2pe_r1_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r1_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR1_0\033[0m -> \033[97mvertex_mm2pe_r1[2]      \033[0m %h", vertex_mm2pe_r1_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r1_3__rst__q1 <= vertex_mm2pe_r1_3__rst__q0;
    vertex_mm2pe_r1_3__rst__q2 <= vertex_mm2pe_r1_3__rst__q1;
  end

  assign vertex_mm2pe_r1_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r1_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r1[3]\033[0m -> \033[90mVertexRouterR2_0        \033[0m %h", vertex_mm2pe_r1_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r1_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR1_0\033[0m -> \033[97mvertex_mm2pe_r1[3]      \033[0m %h", vertex_mm2pe_r1_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r2_0__rst__q1 <= vertex_mm2pe_r2_0__rst__q0;
    vertex_mm2pe_r2_0__rst__q2 <= vertex_mm2pe_r2_0__rst__q1;
  end

  assign vertex_mm2pe_r2_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r2_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r2[0]\033[0m -> \033[90mProcElem_4              \033[0m %h", vertex_mm2pe_r2_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r2_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR2_0\033[0m -> \033[97mvertex_mm2pe_r2[0]      \033[0m %h", vertex_mm2pe_r2_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r2_1__rst__q1 <= vertex_mm2pe_r2_1__rst__q0;
    vertex_mm2pe_r2_1__rst__q2 <= vertex_mm2pe_r2_1__rst__q1;
  end

  assign vertex_mm2pe_r2_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r2_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r2[1]\033[0m -> \033[90mProcElem_5              \033[0m %h", vertex_mm2pe_r2_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r2_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR2_0\033[0m -> \033[97mvertex_mm2pe_r2[1]      \033[0m %h", vertex_mm2pe_r2_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r2_2__rst__q1 <= vertex_mm2pe_r2_2__rst__q0;
    vertex_mm2pe_r2_2__rst__q2 <= vertex_mm2pe_r2_2__rst__q1;
  end

  assign vertex_mm2pe_r2_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r2_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r2[2]\033[0m -> \033[90mProcElem_6              \033[0m %h", vertex_mm2pe_r2_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r2_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR2_0\033[0m -> \033[97mvertex_mm2pe_r2[2]      \033[0m %h", vertex_mm2pe_r2_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_mm2pe_r2_3__rst__q1 <= vertex_mm2pe_r2_3__rst__q0;
    vertex_mm2pe_r2_3__rst__q2 <= vertex_mm2pe_r2_3__rst__q1;
  end

  assign vertex_mm2pe_r2_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r2_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_mm2pe_r2[3]\033[0m -> \033[90mProcElem_7              \033[0m %h", vertex_mm2pe_r2_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_mm2pe_r2_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR2_0\033[0m -> \033[97mvertex_mm2pe_r2[3]      \033[0m %h", vertex_mm2pe_r2_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r0_0__rst__q1 <= vertex_pe2mm_r0_0__rst__q0;
    vertex_pe2mm_r0_0__rst__q2 <= vertex_pe2mm_r0_0__rst__q1;
  end

  assign vertex_pe2mm_r0_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r0_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r0[0]\033[0m -> \033[90mVertexMem_0             \033[0m %h", vertex_pe2mm_r0_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r0_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_0\033[0m -> \033[97mvertex_pe2mm_r0[0]      \033[0m %h", vertex_pe2mm_r0_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r0_1__rst__q1 <= vertex_pe2mm_r0_1__rst__q0;
    vertex_pe2mm_r0_1__rst__q2 <= vertex_pe2mm_r0_1__rst__q1;
  end

  assign vertex_pe2mm_r0_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r0_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r0[1]\033[0m -> \033[90mVertexMem_0             \033[0m %h", vertex_pe2mm_r0_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r0_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR1_0\033[0m -> \033[97mvertex_pe2mm_r0[1]      \033[0m %h", vertex_pe2mm_r0_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r1_0__rst__q1 <= vertex_pe2mm_r1_0__rst__q0;
    vertex_pe2mm_r1_0__rst__q2 <= vertex_pe2mm_r1_0__rst__q1;
  end

  assign vertex_pe2mm_r1_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r1_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r1[0]\033[0m -> \033[90mVertexRouterR1_0        \033[0m %h", vertex_pe2mm_r1_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r1_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_1\033[0m -> \033[97mvertex_pe2mm_r1[0]      \033[0m %h", vertex_pe2mm_r1_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r1_1__rst__q1 <= vertex_pe2mm_r1_1__rst__q0;
    vertex_pe2mm_r1_1__rst__q2 <= vertex_pe2mm_r1_1__rst__q1;
  end

  assign vertex_pe2mm_r1_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r1_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r1[1]\033[0m -> \033[90mVertexRouterR1_0        \033[0m %h", vertex_pe2mm_r1_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r1_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_2\033[0m -> \033[97mvertex_pe2mm_r1[1]      \033[0m %h", vertex_pe2mm_r1_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r1_2__rst__q1 <= vertex_pe2mm_r1_2__rst__q0;
    vertex_pe2mm_r1_2__rst__q2 <= vertex_pe2mm_r1_2__rst__q1;
  end

  assign vertex_pe2mm_r1_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r1_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r1[2]\033[0m -> \033[90mVertexRouterR1_0        \033[0m %h", vertex_pe2mm_r1_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r1_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_3\033[0m -> \033[97mvertex_pe2mm_r1[2]      \033[0m %h", vertex_pe2mm_r1_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r1_3__rst__q1 <= vertex_pe2mm_r1_3__rst__q0;
    vertex_pe2mm_r1_3__rst__q2 <= vertex_pe2mm_r1_3__rst__q1;
  end

  assign vertex_pe2mm_r1_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r1_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r1[3]\033[0m -> \033[90mVertexRouterR1_0        \033[0m %h", vertex_pe2mm_r1_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r1_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR2_0\033[0m -> \033[97mvertex_pe2mm_r1[3]      \033[0m %h", vertex_pe2mm_r1_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r2_0__rst__q1 <= vertex_pe2mm_r2_0__rst__q0;
    vertex_pe2mm_r2_0__rst__q2 <= vertex_pe2mm_r2_0__rst__q1;
  end

  assign vertex_pe2mm_r2_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r2_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r2[0]\033[0m -> \033[90mVertexRouterR2_0        \033[0m %h", vertex_pe2mm_r2_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r2_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_4\033[0m -> \033[97mvertex_pe2mm_r2[0]      \033[0m %h", vertex_pe2mm_r2_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r2_1__rst__q1 <= vertex_pe2mm_r2_1__rst__q0;
    vertex_pe2mm_r2_1__rst__q2 <= vertex_pe2mm_r2_1__rst__q1;
  end

  assign vertex_pe2mm_r2_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r2_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r2[1]\033[0m -> \033[90mVertexRouterR2_0        \033[0m %h", vertex_pe2mm_r2_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r2_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_5\033[0m -> \033[97mvertex_pe2mm_r2[1]      \033[0m %h", vertex_pe2mm_r2_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r2_2__rst__q1 <= vertex_pe2mm_r2_2__rst__q0;
    vertex_pe2mm_r2_2__rst__q2 <= vertex_pe2mm_r2_2__rst__q1;
  end

  assign vertex_pe2mm_r2_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r2_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r2[2]\033[0m -> \033[90mVertexRouterR2_0        \033[0m %h", vertex_pe2mm_r2_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r2_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_6\033[0m -> \033[97mvertex_pe2mm_r2[2]      \033[0m %h", vertex_pe2mm_r2_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_pe2mm_r2_3__rst__q1 <= vertex_pe2mm_r2_3__rst__q0;
    vertex_pe2mm_r2_3__rst__q2 <= vertex_pe2mm_r2_3__rst__q1;
  end

  assign vertex_pe2mm_r2_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r2_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m      vertex_pe2mm_r2[3]\033[0m -> \033[90mVertexRouterR2_0        \033[0m %h", vertex_pe2mm_r2_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_pe2mm_r2_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_7\033[0m -> \033[97mvertex_pe2mm_r2[3]      \033[0m %h", vertex_pe2mm_r2_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r0_0__rst__q1 <= vertex_req_r0_0__rst__q0;
    vertex_req_r0_0__rst__q2 <= vertex_req_r0_0__rst__q1;
  end

  assign vertex_req_r0_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r0_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r0[0]\033[0m -> \033[90mVertexMem_0             \033[0m %h", vertex_req_r0_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r0_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_0\033[0m -> \033[97mvertex_req_r0[0]        \033[0m %h", vertex_req_r0_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r0_1__rst__q1 <= vertex_req_r0_1__rst__q0;
    vertex_req_r0_1__rst__q2 <= vertex_req_r0_1__rst__q1;
  end

  assign vertex_req_r0_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r0_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r0[1]\033[0m -> \033[90mVertexMem_0             \033[0m %h", vertex_req_r0_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r0_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR1_0\033[0m -> \033[97mvertex_req_r0[1]        \033[0m %h", vertex_req_r0_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r1_0__rst__q1 <= vertex_req_r1_0__rst__q0;
    vertex_req_r1_0__rst__q2 <= vertex_req_r1_0__rst__q1;
  end

  assign vertex_req_r1_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r1_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r1[0]\033[0m -> \033[90mVertexRouterR1_0        \033[0m %h", vertex_req_r1_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r1_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_1\033[0m -> \033[97mvertex_req_r1[0]        \033[0m %h", vertex_req_r1_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r1_1__rst__q1 <= vertex_req_r1_1__rst__q0;
    vertex_req_r1_1__rst__q2 <= vertex_req_r1_1__rst__q1;
  end

  assign vertex_req_r1_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r1_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r1[1]\033[0m -> \033[90mVertexRouterR1_0        \033[0m %h", vertex_req_r1_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r1_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_2\033[0m -> \033[97mvertex_req_r1[1]        \033[0m %h", vertex_req_r1_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r1_2__rst__q1 <= vertex_req_r1_2__rst__q0;
    vertex_req_r1_2__rst__q2 <= vertex_req_r1_2__rst__q1;
  end

  assign vertex_req_r1_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r1_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r1[2]\033[0m -> \033[90mVertexRouterR1_0        \033[0m %h", vertex_req_r1_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r1_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_3\033[0m -> \033[97mvertex_req_r1[2]        \033[0m %h", vertex_req_r1_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r1_3__rst__q1 <= vertex_req_r1_3__rst__q0;
    vertex_req_r1_3__rst__q2 <= vertex_req_r1_3__rst__q1;
  end

  assign vertex_req_r1_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r1_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r1[3]\033[0m -> \033[90mVertexRouterR1_0        \033[0m %h", vertex_req_r1_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r1_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m        VertexRouterR2_0\033[0m -> \033[97mvertex_req_r1[3]        \033[0m %h", vertex_req_r1_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r2_0__rst__q1 <= vertex_req_r2_0__rst__q0;
    vertex_req_r2_0__rst__q2 <= vertex_req_r2_0__rst__q1;
  end

  assign vertex_req_r2_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r2_0__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r2[0]\033[0m -> \033[90mVertexRouterR2_0        \033[0m %h", vertex_req_r2_0__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r2_0__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_4\033[0m -> \033[97mvertex_req_r2[0]        \033[0m %h", vertex_req_r2_0__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r2_1__rst__q1 <= vertex_req_r2_1__rst__q0;
    vertex_req_r2_1__rst__q2 <= vertex_req_r2_1__rst__q1;
  end

  assign vertex_req_r2_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r2_1__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r2[1]\033[0m -> \033[90mVertexRouterR2_0        \033[0m %h", vertex_req_r2_1__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r2_1__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_5\033[0m -> \033[97mvertex_req_r2[1]        \033[0m %h", vertex_req_r2_1__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r2_2__rst__q1 <= vertex_req_r2_2__rst__q0;
    vertex_req_r2_2__rst__q2 <= vertex_req_r2_2__rst__q1;
  end

  assign vertex_req_r2_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r2_2__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r2[2]\033[0m -> \033[90mVertexRouterR2_0        \033[0m %h", vertex_req_r2_2__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r2_2__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_6\033[0m -> \033[97mvertex_req_r2[2]        \033[0m %h", vertex_req_r2_2__din);
    end 
  end


  always @(posedge ap_clk) begin
    vertex_req_r2_3__rst__q1 <= vertex_req_r2_3__rst__q0;
    vertex_req_r2_3__rst__q2 <= vertex_req_r2_3__rst__q1;
  end

  assign vertex_req_r2_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(vertex_req_r2_3__read == 1'b1) begin
      $display("DEBUG: R: \033[97m        vertex_req_r2[3]\033[0m -> \033[90mVertexRouterR2_0        \033[0m %h", vertex_req_r2_3__dout);
    end 
  end


  always @(posedge ap_clk) begin
    if(vertex_req_r2_3__write == 1'b1) begin
      $display("DEBUG: W: \033[90m              ProcElem_7\033[0m -> \033[97mvertex_req_r2[3]        \033[0m %h", vertex_req_r2_3__din);
    end 
  end


  always @(posedge ap_clk) begin
    metadata__q1 <= metadata__q0;
    metadata__q2 <= metadata__q1;
  end

  assign metadata__q0 = metadata;

  always @(posedge ap_clk) begin
    Control_0___num_partitions__q1 <= Control_0___num_partitions__q0;
    Control_0___num_partitions__q2 <= Control_0___num_partitions__q1;
  end

  assign Control_0___num_partitions__q0 = num_partitions;

  always @(posedge ap_clk) begin
    Control_0__ap_rst_n__q1 <= Control_0__ap_rst_n__q0;
    Control_0__ap_rst_n__q2 <= Control_0__ap_rst_n__q1;
  end

  assign Control_0__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    Control_0__is_done__q1 <= Control_0__is_done__q0;
    Control_0__is_done__q2 <= Control_0__is_done__q1;
  end

  assign Control_0__is_done__q0 = (Control_0__state == 2'b10);

  always @(posedge ap_clk) begin
    Control_0__ap_start_global__q1 <= Control_0__ap_start_global__q0;
    Control_0__ap_start_global__q2 <= Control_0__ap_start_global__q1;
  end

  assign Control_0__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    Control_0__ap_done_global__q1 <= Control_0__ap_done_global__q0;
    Control_0__ap_done_global__q2 <= Control_0__ap_done_global__q1;
  end

  assign Control_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~Control_0__ap_rst_n__q2) begin
      Control_0__state <= 2'b00;
    end else begin
      if(Control_0__state == 2'b00) begin
        if(Control_0__ap_start_global__q2) begin
          Control_0__state <= 2'b01;
        end 
      end 
      if(Control_0__state == 2'b01) begin
        if(Control_0__ap_ready) begin
          if(Control_0__ap_done) begin
            Control_0__state <= 2'b10;
          end else begin
            Control_0__state <= 2'b11;
          end
        end 
      end 
      if(Control_0__state == 2'b11) begin
        if(Control_0__ap_done) begin
          Control_0__state <= 2'b10;
        end 
      end 
      if(Control_0__state == 2'b10) begin
        if(Control_0__ap_done_global__q2) begin
          Control_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign Control_0__ap_start = (Control_0__state == 2'b01);

  always @(posedge ap_clk) begin
    edges_0__q1 <= edges_0__q0;
    edges_0__q2 <= edges_0__q1;
  end

  assign edges_0__q0 = edges_0;

  always @(posedge ap_clk) begin
    EdgeMem_0__ap_rst_n__q1 <= EdgeMem_0__ap_rst_n__q0;
    EdgeMem_0__ap_rst_n__q2 <= EdgeMem_0__ap_rst_n__q1;
  end

  assign EdgeMem_0__ap_rst_n__q0 = ap_rst_n;
  assign EdgeMem_0__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    edges_1__q1 <= edges_1__q0;
    edges_1__q2 <= edges_1__q1;
  end

  assign edges_1__q0 = edges_1;

  always @(posedge ap_clk) begin
    EdgeMem_1__ap_rst_n__q1 <= EdgeMem_1__ap_rst_n__q0;
    EdgeMem_1__ap_rst_n__q2 <= EdgeMem_1__ap_rst_n__q1;
  end

  assign EdgeMem_1__ap_rst_n__q0 = ap_rst_n;
  assign EdgeMem_1__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    edges_2__q1 <= edges_2__q0;
    edges_2__q2 <= edges_2__q1;
  end

  assign edges_2__q0 = edges_2;

  always @(posedge ap_clk) begin
    EdgeMem_2__ap_rst_n__q1 <= EdgeMem_2__ap_rst_n__q0;
    EdgeMem_2__ap_rst_n__q2 <= EdgeMem_2__ap_rst_n__q1;
  end

  assign EdgeMem_2__ap_rst_n__q0 = ap_rst_n;
  assign EdgeMem_2__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    edges_3__q1 <= edges_3__q0;
    edges_3__q2 <= edges_3__q1;
  end

  assign edges_3__q0 = edges_3;

  always @(posedge ap_clk) begin
    EdgeMem_3__ap_rst_n__q1 <= EdgeMem_3__ap_rst_n__q0;
    EdgeMem_3__ap_rst_n__q2 <= EdgeMem_3__ap_rst_n__q1;
  end

  assign EdgeMem_3__ap_rst_n__q0 = ap_rst_n;
  assign EdgeMem_3__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    edges_4__q1 <= edges_4__q0;
    edges_4__q2 <= edges_4__q1;
  end

  assign edges_4__q0 = edges_4;

  always @(posedge ap_clk) begin
    EdgeMem_4__ap_rst_n__q1 <= EdgeMem_4__ap_rst_n__q0;
    EdgeMem_4__ap_rst_n__q2 <= EdgeMem_4__ap_rst_n__q1;
  end

  assign EdgeMem_4__ap_rst_n__q0 = ap_rst_n;
  assign EdgeMem_4__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    edges_5__q1 <= edges_5__q0;
    edges_5__q2 <= edges_5__q1;
  end

  assign edges_5__q0 = edges_5;

  always @(posedge ap_clk) begin
    EdgeMem_5__ap_rst_n__q1 <= EdgeMem_5__ap_rst_n__q0;
    EdgeMem_5__ap_rst_n__q2 <= EdgeMem_5__ap_rst_n__q1;
  end

  assign EdgeMem_5__ap_rst_n__q0 = ap_rst_n;
  assign EdgeMem_5__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    edges_6__q1 <= edges_6__q0;
    edges_6__q2 <= edges_6__q1;
  end

  assign edges_6__q0 = edges_6;

  always @(posedge ap_clk) begin
    EdgeMem_6__ap_rst_n__q1 <= EdgeMem_6__ap_rst_n__q0;
    EdgeMem_6__ap_rst_n__q2 <= EdgeMem_6__ap_rst_n__q1;
  end

  assign EdgeMem_6__ap_rst_n__q0 = ap_rst_n;
  assign EdgeMem_6__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    edges_7__q1 <= edges_7__q0;
    edges_7__q2 <= edges_7__q1;
  end

  assign edges_7__q0 = edges_7;

  always @(posedge ap_clk) begin
    EdgeMem_7__ap_rst_n__q1 <= EdgeMem_7__ap_rst_n__q0;
    EdgeMem_7__ap_rst_n__q2 <= EdgeMem_7__ap_rst_n__q1;
  end

  assign EdgeMem_7__ap_rst_n__q0 = ap_rst_n;
  assign EdgeMem_7__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    ProcElem_0__ap_rst_n__q1 <= ProcElem_0__ap_rst_n__q0;
    ProcElem_0__ap_rst_n__q2 <= ProcElem_0__ap_rst_n__q1;
  end

  assign ProcElem_0__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    ProcElem_0__is_done__q1 <= ProcElem_0__is_done__q0;
    ProcElem_0__is_done__q2 <= ProcElem_0__is_done__q1;
  end

  assign ProcElem_0__is_done__q0 = (ProcElem_0__state == 2'b10);

  always @(posedge ap_clk) begin
    ProcElem_0__ap_start_global__q1 <= ProcElem_0__ap_start_global__q0;
    ProcElem_0__ap_start_global__q2 <= ProcElem_0__ap_start_global__q1;
  end

  assign ProcElem_0__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    ProcElem_0__ap_done_global__q1 <= ProcElem_0__ap_done_global__q0;
    ProcElem_0__ap_done_global__q2 <= ProcElem_0__ap_done_global__q1;
  end

  assign ProcElem_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ProcElem_0__ap_rst_n__q2) begin
      ProcElem_0__state <= 2'b00;
    end else begin
      if(ProcElem_0__state == 2'b00) begin
        if(ProcElem_0__ap_start_global__q2) begin
          ProcElem_0__state <= 2'b01;
        end 
      end 
      if(ProcElem_0__state == 2'b01) begin
        if(ProcElem_0__ap_ready) begin
          if(ProcElem_0__ap_done) begin
            ProcElem_0__state <= 2'b10;
          end else begin
            ProcElem_0__state <= 2'b11;
          end
        end 
      end 
      if(ProcElem_0__state == 2'b11) begin
        if(ProcElem_0__ap_done) begin
          ProcElem_0__state <= 2'b10;
        end 
      end 
      if(ProcElem_0__state == 2'b10) begin
        if(ProcElem_0__ap_done_global__q2) begin
          ProcElem_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign ProcElem_0__ap_start = (ProcElem_0__state == 2'b01);

  always @(posedge ap_clk) begin
    ProcElem_1__ap_rst_n__q1 <= ProcElem_1__ap_rst_n__q0;
    ProcElem_1__ap_rst_n__q2 <= ProcElem_1__ap_rst_n__q1;
  end

  assign ProcElem_1__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    ProcElem_1__is_done__q1 <= ProcElem_1__is_done__q0;
    ProcElem_1__is_done__q2 <= ProcElem_1__is_done__q1;
  end

  assign ProcElem_1__is_done__q0 = (ProcElem_1__state == 2'b10);

  always @(posedge ap_clk) begin
    ProcElem_1__ap_start_global__q1 <= ProcElem_1__ap_start_global__q0;
    ProcElem_1__ap_start_global__q2 <= ProcElem_1__ap_start_global__q1;
  end

  assign ProcElem_1__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    ProcElem_1__ap_done_global__q1 <= ProcElem_1__ap_done_global__q0;
    ProcElem_1__ap_done_global__q2 <= ProcElem_1__ap_done_global__q1;
  end

  assign ProcElem_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ProcElem_1__ap_rst_n__q2) begin
      ProcElem_1__state <= 2'b00;
    end else begin
      if(ProcElem_1__state == 2'b00) begin
        if(ProcElem_1__ap_start_global__q2) begin
          ProcElem_1__state <= 2'b01;
        end 
      end 
      if(ProcElem_1__state == 2'b01) begin
        if(ProcElem_1__ap_ready) begin
          if(ProcElem_1__ap_done) begin
            ProcElem_1__state <= 2'b10;
          end else begin
            ProcElem_1__state <= 2'b11;
          end
        end 
      end 
      if(ProcElem_1__state == 2'b11) begin
        if(ProcElem_1__ap_done) begin
          ProcElem_1__state <= 2'b10;
        end 
      end 
      if(ProcElem_1__state == 2'b10) begin
        if(ProcElem_1__ap_done_global__q2) begin
          ProcElem_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign ProcElem_1__ap_start = (ProcElem_1__state == 2'b01);

  always @(posedge ap_clk) begin
    ProcElem_2__ap_rst_n__q1 <= ProcElem_2__ap_rst_n__q0;
    ProcElem_2__ap_rst_n__q2 <= ProcElem_2__ap_rst_n__q1;
  end

  assign ProcElem_2__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    ProcElem_2__is_done__q1 <= ProcElem_2__is_done__q0;
    ProcElem_2__is_done__q2 <= ProcElem_2__is_done__q1;
  end

  assign ProcElem_2__is_done__q0 = (ProcElem_2__state == 2'b10);

  always @(posedge ap_clk) begin
    ProcElem_2__ap_start_global__q1 <= ProcElem_2__ap_start_global__q0;
    ProcElem_2__ap_start_global__q2 <= ProcElem_2__ap_start_global__q1;
  end

  assign ProcElem_2__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    ProcElem_2__ap_done_global__q1 <= ProcElem_2__ap_done_global__q0;
    ProcElem_2__ap_done_global__q2 <= ProcElem_2__ap_done_global__q1;
  end

  assign ProcElem_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ProcElem_2__ap_rst_n__q2) begin
      ProcElem_2__state <= 2'b00;
    end else begin
      if(ProcElem_2__state == 2'b00) begin
        if(ProcElem_2__ap_start_global__q2) begin
          ProcElem_2__state <= 2'b01;
        end 
      end 
      if(ProcElem_2__state == 2'b01) begin
        if(ProcElem_2__ap_ready) begin
          if(ProcElem_2__ap_done) begin
            ProcElem_2__state <= 2'b10;
          end else begin
            ProcElem_2__state <= 2'b11;
          end
        end 
      end 
      if(ProcElem_2__state == 2'b11) begin
        if(ProcElem_2__ap_done) begin
          ProcElem_2__state <= 2'b10;
        end 
      end 
      if(ProcElem_2__state == 2'b10) begin
        if(ProcElem_2__ap_done_global__q2) begin
          ProcElem_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign ProcElem_2__ap_start = (ProcElem_2__state == 2'b01);

  always @(posedge ap_clk) begin
    ProcElem_3__ap_rst_n__q1 <= ProcElem_3__ap_rst_n__q0;
    ProcElem_3__ap_rst_n__q2 <= ProcElem_3__ap_rst_n__q1;
  end

  assign ProcElem_3__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    ProcElem_3__is_done__q1 <= ProcElem_3__is_done__q0;
    ProcElem_3__is_done__q2 <= ProcElem_3__is_done__q1;
  end

  assign ProcElem_3__is_done__q0 = (ProcElem_3__state == 2'b10);

  always @(posedge ap_clk) begin
    ProcElem_3__ap_start_global__q1 <= ProcElem_3__ap_start_global__q0;
    ProcElem_3__ap_start_global__q2 <= ProcElem_3__ap_start_global__q1;
  end

  assign ProcElem_3__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    ProcElem_3__ap_done_global__q1 <= ProcElem_3__ap_done_global__q0;
    ProcElem_3__ap_done_global__q2 <= ProcElem_3__ap_done_global__q1;
  end

  assign ProcElem_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ProcElem_3__ap_rst_n__q2) begin
      ProcElem_3__state <= 2'b00;
    end else begin
      if(ProcElem_3__state == 2'b00) begin
        if(ProcElem_3__ap_start_global__q2) begin
          ProcElem_3__state <= 2'b01;
        end 
      end 
      if(ProcElem_3__state == 2'b01) begin
        if(ProcElem_3__ap_ready) begin
          if(ProcElem_3__ap_done) begin
            ProcElem_3__state <= 2'b10;
          end else begin
            ProcElem_3__state <= 2'b11;
          end
        end 
      end 
      if(ProcElem_3__state == 2'b11) begin
        if(ProcElem_3__ap_done) begin
          ProcElem_3__state <= 2'b10;
        end 
      end 
      if(ProcElem_3__state == 2'b10) begin
        if(ProcElem_3__ap_done_global__q2) begin
          ProcElem_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign ProcElem_3__ap_start = (ProcElem_3__state == 2'b01);

  always @(posedge ap_clk) begin
    ProcElem_4__ap_rst_n__q1 <= ProcElem_4__ap_rst_n__q0;
    ProcElem_4__ap_rst_n__q2 <= ProcElem_4__ap_rst_n__q1;
  end

  assign ProcElem_4__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    ProcElem_4__is_done__q1 <= ProcElem_4__is_done__q0;
    ProcElem_4__is_done__q2 <= ProcElem_4__is_done__q1;
  end

  assign ProcElem_4__is_done__q0 = (ProcElem_4__state == 2'b10);

  always @(posedge ap_clk) begin
    ProcElem_4__ap_start_global__q1 <= ProcElem_4__ap_start_global__q0;
    ProcElem_4__ap_start_global__q2 <= ProcElem_4__ap_start_global__q1;
  end

  assign ProcElem_4__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    ProcElem_4__ap_done_global__q1 <= ProcElem_4__ap_done_global__q0;
    ProcElem_4__ap_done_global__q2 <= ProcElem_4__ap_done_global__q1;
  end

  assign ProcElem_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ProcElem_4__ap_rst_n__q2) begin
      ProcElem_4__state <= 2'b00;
    end else begin
      if(ProcElem_4__state == 2'b00) begin
        if(ProcElem_4__ap_start_global__q2) begin
          ProcElem_4__state <= 2'b01;
        end 
      end 
      if(ProcElem_4__state == 2'b01) begin
        if(ProcElem_4__ap_ready) begin
          if(ProcElem_4__ap_done) begin
            ProcElem_4__state <= 2'b10;
          end else begin
            ProcElem_4__state <= 2'b11;
          end
        end 
      end 
      if(ProcElem_4__state == 2'b11) begin
        if(ProcElem_4__ap_done) begin
          ProcElem_4__state <= 2'b10;
        end 
      end 
      if(ProcElem_4__state == 2'b10) begin
        if(ProcElem_4__ap_done_global__q2) begin
          ProcElem_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign ProcElem_4__ap_start = (ProcElem_4__state == 2'b01);

  always @(posedge ap_clk) begin
    ProcElem_5__ap_rst_n__q1 <= ProcElem_5__ap_rst_n__q0;
    ProcElem_5__ap_rst_n__q2 <= ProcElem_5__ap_rst_n__q1;
  end

  assign ProcElem_5__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    ProcElem_5__is_done__q1 <= ProcElem_5__is_done__q0;
    ProcElem_5__is_done__q2 <= ProcElem_5__is_done__q1;
  end

  assign ProcElem_5__is_done__q0 = (ProcElem_5__state == 2'b10);

  always @(posedge ap_clk) begin
    ProcElem_5__ap_start_global__q1 <= ProcElem_5__ap_start_global__q0;
    ProcElem_5__ap_start_global__q2 <= ProcElem_5__ap_start_global__q1;
  end

  assign ProcElem_5__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    ProcElem_5__ap_done_global__q1 <= ProcElem_5__ap_done_global__q0;
    ProcElem_5__ap_done_global__q2 <= ProcElem_5__ap_done_global__q1;
  end

  assign ProcElem_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ProcElem_5__ap_rst_n__q2) begin
      ProcElem_5__state <= 2'b00;
    end else begin
      if(ProcElem_5__state == 2'b00) begin
        if(ProcElem_5__ap_start_global__q2) begin
          ProcElem_5__state <= 2'b01;
        end 
      end 
      if(ProcElem_5__state == 2'b01) begin
        if(ProcElem_5__ap_ready) begin
          if(ProcElem_5__ap_done) begin
            ProcElem_5__state <= 2'b10;
          end else begin
            ProcElem_5__state <= 2'b11;
          end
        end 
      end 
      if(ProcElem_5__state == 2'b11) begin
        if(ProcElem_5__ap_done) begin
          ProcElem_5__state <= 2'b10;
        end 
      end 
      if(ProcElem_5__state == 2'b10) begin
        if(ProcElem_5__ap_done_global__q2) begin
          ProcElem_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign ProcElem_5__ap_start = (ProcElem_5__state == 2'b01);

  always @(posedge ap_clk) begin
    ProcElem_6__ap_rst_n__q1 <= ProcElem_6__ap_rst_n__q0;
    ProcElem_6__ap_rst_n__q2 <= ProcElem_6__ap_rst_n__q1;
  end

  assign ProcElem_6__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    ProcElem_6__is_done__q1 <= ProcElem_6__is_done__q0;
    ProcElem_6__is_done__q2 <= ProcElem_6__is_done__q1;
  end

  assign ProcElem_6__is_done__q0 = (ProcElem_6__state == 2'b10);

  always @(posedge ap_clk) begin
    ProcElem_6__ap_start_global__q1 <= ProcElem_6__ap_start_global__q0;
    ProcElem_6__ap_start_global__q2 <= ProcElem_6__ap_start_global__q1;
  end

  assign ProcElem_6__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    ProcElem_6__ap_done_global__q1 <= ProcElem_6__ap_done_global__q0;
    ProcElem_6__ap_done_global__q2 <= ProcElem_6__ap_done_global__q1;
  end

  assign ProcElem_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ProcElem_6__ap_rst_n__q2) begin
      ProcElem_6__state <= 2'b00;
    end else begin
      if(ProcElem_6__state == 2'b00) begin
        if(ProcElem_6__ap_start_global__q2) begin
          ProcElem_6__state <= 2'b01;
        end 
      end 
      if(ProcElem_6__state == 2'b01) begin
        if(ProcElem_6__ap_ready) begin
          if(ProcElem_6__ap_done) begin
            ProcElem_6__state <= 2'b10;
          end else begin
            ProcElem_6__state <= 2'b11;
          end
        end 
      end 
      if(ProcElem_6__state == 2'b11) begin
        if(ProcElem_6__ap_done) begin
          ProcElem_6__state <= 2'b10;
        end 
      end 
      if(ProcElem_6__state == 2'b10) begin
        if(ProcElem_6__ap_done_global__q2) begin
          ProcElem_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign ProcElem_6__ap_start = (ProcElem_6__state == 2'b01);

  always @(posedge ap_clk) begin
    ProcElem_7__ap_rst_n__q1 <= ProcElem_7__ap_rst_n__q0;
    ProcElem_7__ap_rst_n__q2 <= ProcElem_7__ap_rst_n__q1;
  end

  assign ProcElem_7__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    ProcElem_7__is_done__q1 <= ProcElem_7__is_done__q0;
    ProcElem_7__is_done__q2 <= ProcElem_7__is_done__q1;
  end

  assign ProcElem_7__is_done__q0 = (ProcElem_7__state == 2'b10);

  always @(posedge ap_clk) begin
    ProcElem_7__ap_start_global__q1 <= ProcElem_7__ap_start_global__q0;
    ProcElem_7__ap_start_global__q2 <= ProcElem_7__ap_start_global__q1;
  end

  assign ProcElem_7__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    ProcElem_7__ap_done_global__q1 <= ProcElem_7__ap_done_global__q0;
    ProcElem_7__ap_done_global__q2 <= ProcElem_7__ap_done_global__q1;
  end

  assign ProcElem_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ProcElem_7__ap_rst_n__q2) begin
      ProcElem_7__state <= 2'b00;
    end else begin
      if(ProcElem_7__state == 2'b00) begin
        if(ProcElem_7__ap_start_global__q2) begin
          ProcElem_7__state <= 2'b01;
        end 
      end 
      if(ProcElem_7__state == 2'b01) begin
        if(ProcElem_7__ap_ready) begin
          if(ProcElem_7__ap_done) begin
            ProcElem_7__state <= 2'b10;
          end else begin
            ProcElem_7__state <= 2'b11;
          end
        end 
      end 
      if(ProcElem_7__state == 2'b11) begin
        if(ProcElem_7__ap_done) begin
          ProcElem_7__state <= 2'b10;
        end 
      end 
      if(ProcElem_7__state == 2'b10) begin
        if(ProcElem_7__ap_done_global__q2) begin
          ProcElem_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign ProcElem_7__ap_start = (ProcElem_7__state == 2'b01);

  always @(posedge ap_clk) begin
    UpdateHandler_0___num_partitions__q1 <= UpdateHandler_0___num_partitions__q0;
    UpdateHandler_0___num_partitions__q2 <= UpdateHandler_0___num_partitions__q1;
  end

  assign UpdateHandler_0___num_partitions__q0 = num_partitions;

  always @(posedge ap_clk) begin
    UpdateHandler_0__ap_rst_n__q1 <= UpdateHandler_0__ap_rst_n__q0;
    UpdateHandler_0__ap_rst_n__q2 <= UpdateHandler_0__ap_rst_n__q1;
  end

  assign UpdateHandler_0__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    UpdateHandler_0__is_done__q1 <= UpdateHandler_0__is_done__q0;
    UpdateHandler_0__is_done__q2 <= UpdateHandler_0__is_done__q1;
  end

  assign UpdateHandler_0__is_done__q0 = (UpdateHandler_0__state == 2'b10);

  always @(posedge ap_clk) begin
    UpdateHandler_0__ap_start_global__q1 <= UpdateHandler_0__ap_start_global__q0;
    UpdateHandler_0__ap_start_global__q2 <= UpdateHandler_0__ap_start_global__q1;
  end

  assign UpdateHandler_0__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    UpdateHandler_0__ap_done_global__q1 <= UpdateHandler_0__ap_done_global__q0;
    UpdateHandler_0__ap_done_global__q2 <= UpdateHandler_0__ap_done_global__q1;
  end

  assign UpdateHandler_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~UpdateHandler_0__ap_rst_n__q2) begin
      UpdateHandler_0__state <= 2'b00;
    end else begin
      if(UpdateHandler_0__state == 2'b00) begin
        if(UpdateHandler_0__ap_start_global__q2) begin
          UpdateHandler_0__state <= 2'b01;
        end 
      end 
      if(UpdateHandler_0__state == 2'b01) begin
        if(UpdateHandler_0__ap_ready) begin
          if(UpdateHandler_0__ap_done) begin
            UpdateHandler_0__state <= 2'b10;
          end else begin
            UpdateHandler_0__state <= 2'b11;
          end
        end 
      end 
      if(UpdateHandler_0__state == 2'b11) begin
        if(UpdateHandler_0__ap_done) begin
          UpdateHandler_0__state <= 2'b10;
        end 
      end 
      if(UpdateHandler_0__state == 2'b10) begin
        if(UpdateHandler_0__ap_done_global__q2) begin
          UpdateHandler_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign UpdateHandler_0__ap_start = (UpdateHandler_0__state == 2'b01);

  always @(posedge ap_clk) begin
    UpdateHandler_1___num_partitions__q1 <= UpdateHandler_1___num_partitions__q0;
    UpdateHandler_1___num_partitions__q2 <= UpdateHandler_1___num_partitions__q1;
  end

  assign UpdateHandler_1___num_partitions__q0 = num_partitions;

  always @(posedge ap_clk) begin
    UpdateHandler_1__ap_rst_n__q1 <= UpdateHandler_1__ap_rst_n__q0;
    UpdateHandler_1__ap_rst_n__q2 <= UpdateHandler_1__ap_rst_n__q1;
  end

  assign UpdateHandler_1__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    UpdateHandler_1__is_done__q1 <= UpdateHandler_1__is_done__q0;
    UpdateHandler_1__is_done__q2 <= UpdateHandler_1__is_done__q1;
  end

  assign UpdateHandler_1__is_done__q0 = (UpdateHandler_1__state == 2'b10);

  always @(posedge ap_clk) begin
    UpdateHandler_1__ap_start_global__q1 <= UpdateHandler_1__ap_start_global__q0;
    UpdateHandler_1__ap_start_global__q2 <= UpdateHandler_1__ap_start_global__q1;
  end

  assign UpdateHandler_1__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    UpdateHandler_1__ap_done_global__q1 <= UpdateHandler_1__ap_done_global__q0;
    UpdateHandler_1__ap_done_global__q2 <= UpdateHandler_1__ap_done_global__q1;
  end

  assign UpdateHandler_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~UpdateHandler_1__ap_rst_n__q2) begin
      UpdateHandler_1__state <= 2'b00;
    end else begin
      if(UpdateHandler_1__state == 2'b00) begin
        if(UpdateHandler_1__ap_start_global__q2) begin
          UpdateHandler_1__state <= 2'b01;
        end 
      end 
      if(UpdateHandler_1__state == 2'b01) begin
        if(UpdateHandler_1__ap_ready) begin
          if(UpdateHandler_1__ap_done) begin
            UpdateHandler_1__state <= 2'b10;
          end else begin
            UpdateHandler_1__state <= 2'b11;
          end
        end 
      end 
      if(UpdateHandler_1__state == 2'b11) begin
        if(UpdateHandler_1__ap_done) begin
          UpdateHandler_1__state <= 2'b10;
        end 
      end 
      if(UpdateHandler_1__state == 2'b10) begin
        if(UpdateHandler_1__ap_done_global__q2) begin
          UpdateHandler_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign UpdateHandler_1__ap_start = (UpdateHandler_1__state == 2'b01);

  always @(posedge ap_clk) begin
    UpdateHandler_2___num_partitions__q1 <= UpdateHandler_2___num_partitions__q0;
    UpdateHandler_2___num_partitions__q2 <= UpdateHandler_2___num_partitions__q1;
  end

  assign UpdateHandler_2___num_partitions__q0 = num_partitions;

  always @(posedge ap_clk) begin
    UpdateHandler_2__ap_rst_n__q1 <= UpdateHandler_2__ap_rst_n__q0;
    UpdateHandler_2__ap_rst_n__q2 <= UpdateHandler_2__ap_rst_n__q1;
  end

  assign UpdateHandler_2__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    UpdateHandler_2__is_done__q1 <= UpdateHandler_2__is_done__q0;
    UpdateHandler_2__is_done__q2 <= UpdateHandler_2__is_done__q1;
  end

  assign UpdateHandler_2__is_done__q0 = (UpdateHandler_2__state == 2'b10);

  always @(posedge ap_clk) begin
    UpdateHandler_2__ap_start_global__q1 <= UpdateHandler_2__ap_start_global__q0;
    UpdateHandler_2__ap_start_global__q2 <= UpdateHandler_2__ap_start_global__q1;
  end

  assign UpdateHandler_2__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    UpdateHandler_2__ap_done_global__q1 <= UpdateHandler_2__ap_done_global__q0;
    UpdateHandler_2__ap_done_global__q2 <= UpdateHandler_2__ap_done_global__q1;
  end

  assign UpdateHandler_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~UpdateHandler_2__ap_rst_n__q2) begin
      UpdateHandler_2__state <= 2'b00;
    end else begin
      if(UpdateHandler_2__state == 2'b00) begin
        if(UpdateHandler_2__ap_start_global__q2) begin
          UpdateHandler_2__state <= 2'b01;
        end 
      end 
      if(UpdateHandler_2__state == 2'b01) begin
        if(UpdateHandler_2__ap_ready) begin
          if(UpdateHandler_2__ap_done) begin
            UpdateHandler_2__state <= 2'b10;
          end else begin
            UpdateHandler_2__state <= 2'b11;
          end
        end 
      end 
      if(UpdateHandler_2__state == 2'b11) begin
        if(UpdateHandler_2__ap_done) begin
          UpdateHandler_2__state <= 2'b10;
        end 
      end 
      if(UpdateHandler_2__state == 2'b10) begin
        if(UpdateHandler_2__ap_done_global__q2) begin
          UpdateHandler_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign UpdateHandler_2__ap_start = (UpdateHandler_2__state == 2'b01);

  always @(posedge ap_clk) begin
    UpdateHandler_3___num_partitions__q1 <= UpdateHandler_3___num_partitions__q0;
    UpdateHandler_3___num_partitions__q2 <= UpdateHandler_3___num_partitions__q1;
  end

  assign UpdateHandler_3___num_partitions__q0 = num_partitions;

  always @(posedge ap_clk) begin
    UpdateHandler_3__ap_rst_n__q1 <= UpdateHandler_3__ap_rst_n__q0;
    UpdateHandler_3__ap_rst_n__q2 <= UpdateHandler_3__ap_rst_n__q1;
  end

  assign UpdateHandler_3__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    UpdateHandler_3__is_done__q1 <= UpdateHandler_3__is_done__q0;
    UpdateHandler_3__is_done__q2 <= UpdateHandler_3__is_done__q1;
  end

  assign UpdateHandler_3__is_done__q0 = (UpdateHandler_3__state == 2'b10);

  always @(posedge ap_clk) begin
    UpdateHandler_3__ap_start_global__q1 <= UpdateHandler_3__ap_start_global__q0;
    UpdateHandler_3__ap_start_global__q2 <= UpdateHandler_3__ap_start_global__q1;
  end

  assign UpdateHandler_3__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    UpdateHandler_3__ap_done_global__q1 <= UpdateHandler_3__ap_done_global__q0;
    UpdateHandler_3__ap_done_global__q2 <= UpdateHandler_3__ap_done_global__q1;
  end

  assign UpdateHandler_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~UpdateHandler_3__ap_rst_n__q2) begin
      UpdateHandler_3__state <= 2'b00;
    end else begin
      if(UpdateHandler_3__state == 2'b00) begin
        if(UpdateHandler_3__ap_start_global__q2) begin
          UpdateHandler_3__state <= 2'b01;
        end 
      end 
      if(UpdateHandler_3__state == 2'b01) begin
        if(UpdateHandler_3__ap_ready) begin
          if(UpdateHandler_3__ap_done) begin
            UpdateHandler_3__state <= 2'b10;
          end else begin
            UpdateHandler_3__state <= 2'b11;
          end
        end 
      end 
      if(UpdateHandler_3__state == 2'b11) begin
        if(UpdateHandler_3__ap_done) begin
          UpdateHandler_3__state <= 2'b10;
        end 
      end 
      if(UpdateHandler_3__state == 2'b10) begin
        if(UpdateHandler_3__ap_done_global__q2) begin
          UpdateHandler_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign UpdateHandler_3__ap_start = (UpdateHandler_3__state == 2'b01);

  always @(posedge ap_clk) begin
    UpdateHandler_4___num_partitions__q1 <= UpdateHandler_4___num_partitions__q0;
    UpdateHandler_4___num_partitions__q2 <= UpdateHandler_4___num_partitions__q1;
  end

  assign UpdateHandler_4___num_partitions__q0 = num_partitions;

  always @(posedge ap_clk) begin
    UpdateHandler_4__ap_rst_n__q1 <= UpdateHandler_4__ap_rst_n__q0;
    UpdateHandler_4__ap_rst_n__q2 <= UpdateHandler_4__ap_rst_n__q1;
  end

  assign UpdateHandler_4__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    UpdateHandler_4__is_done__q1 <= UpdateHandler_4__is_done__q0;
    UpdateHandler_4__is_done__q2 <= UpdateHandler_4__is_done__q1;
  end

  assign UpdateHandler_4__is_done__q0 = (UpdateHandler_4__state == 2'b10);

  always @(posedge ap_clk) begin
    UpdateHandler_4__ap_start_global__q1 <= UpdateHandler_4__ap_start_global__q0;
    UpdateHandler_4__ap_start_global__q2 <= UpdateHandler_4__ap_start_global__q1;
  end

  assign UpdateHandler_4__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    UpdateHandler_4__ap_done_global__q1 <= UpdateHandler_4__ap_done_global__q0;
    UpdateHandler_4__ap_done_global__q2 <= UpdateHandler_4__ap_done_global__q1;
  end

  assign UpdateHandler_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~UpdateHandler_4__ap_rst_n__q2) begin
      UpdateHandler_4__state <= 2'b00;
    end else begin
      if(UpdateHandler_4__state == 2'b00) begin
        if(UpdateHandler_4__ap_start_global__q2) begin
          UpdateHandler_4__state <= 2'b01;
        end 
      end 
      if(UpdateHandler_4__state == 2'b01) begin
        if(UpdateHandler_4__ap_ready) begin
          if(UpdateHandler_4__ap_done) begin
            UpdateHandler_4__state <= 2'b10;
          end else begin
            UpdateHandler_4__state <= 2'b11;
          end
        end 
      end 
      if(UpdateHandler_4__state == 2'b11) begin
        if(UpdateHandler_4__ap_done) begin
          UpdateHandler_4__state <= 2'b10;
        end 
      end 
      if(UpdateHandler_4__state == 2'b10) begin
        if(UpdateHandler_4__ap_done_global__q2) begin
          UpdateHandler_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign UpdateHandler_4__ap_start = (UpdateHandler_4__state == 2'b01);

  always @(posedge ap_clk) begin
    UpdateHandler_5___num_partitions__q1 <= UpdateHandler_5___num_partitions__q0;
    UpdateHandler_5___num_partitions__q2 <= UpdateHandler_5___num_partitions__q1;
  end

  assign UpdateHandler_5___num_partitions__q0 = num_partitions;

  always @(posedge ap_clk) begin
    UpdateHandler_5__ap_rst_n__q1 <= UpdateHandler_5__ap_rst_n__q0;
    UpdateHandler_5__ap_rst_n__q2 <= UpdateHandler_5__ap_rst_n__q1;
  end

  assign UpdateHandler_5__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    UpdateHandler_5__is_done__q1 <= UpdateHandler_5__is_done__q0;
    UpdateHandler_5__is_done__q2 <= UpdateHandler_5__is_done__q1;
  end

  assign UpdateHandler_5__is_done__q0 = (UpdateHandler_5__state == 2'b10);

  always @(posedge ap_clk) begin
    UpdateHandler_5__ap_start_global__q1 <= UpdateHandler_5__ap_start_global__q0;
    UpdateHandler_5__ap_start_global__q2 <= UpdateHandler_5__ap_start_global__q1;
  end

  assign UpdateHandler_5__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    UpdateHandler_5__ap_done_global__q1 <= UpdateHandler_5__ap_done_global__q0;
    UpdateHandler_5__ap_done_global__q2 <= UpdateHandler_5__ap_done_global__q1;
  end

  assign UpdateHandler_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~UpdateHandler_5__ap_rst_n__q2) begin
      UpdateHandler_5__state <= 2'b00;
    end else begin
      if(UpdateHandler_5__state == 2'b00) begin
        if(UpdateHandler_5__ap_start_global__q2) begin
          UpdateHandler_5__state <= 2'b01;
        end 
      end 
      if(UpdateHandler_5__state == 2'b01) begin
        if(UpdateHandler_5__ap_ready) begin
          if(UpdateHandler_5__ap_done) begin
            UpdateHandler_5__state <= 2'b10;
          end else begin
            UpdateHandler_5__state <= 2'b11;
          end
        end 
      end 
      if(UpdateHandler_5__state == 2'b11) begin
        if(UpdateHandler_5__ap_done) begin
          UpdateHandler_5__state <= 2'b10;
        end 
      end 
      if(UpdateHandler_5__state == 2'b10) begin
        if(UpdateHandler_5__ap_done_global__q2) begin
          UpdateHandler_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign UpdateHandler_5__ap_start = (UpdateHandler_5__state == 2'b01);

  always @(posedge ap_clk) begin
    UpdateHandler_6___num_partitions__q1 <= UpdateHandler_6___num_partitions__q0;
    UpdateHandler_6___num_partitions__q2 <= UpdateHandler_6___num_partitions__q1;
  end

  assign UpdateHandler_6___num_partitions__q0 = num_partitions;

  always @(posedge ap_clk) begin
    UpdateHandler_6__ap_rst_n__q1 <= UpdateHandler_6__ap_rst_n__q0;
    UpdateHandler_6__ap_rst_n__q2 <= UpdateHandler_6__ap_rst_n__q1;
  end

  assign UpdateHandler_6__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    UpdateHandler_6__is_done__q1 <= UpdateHandler_6__is_done__q0;
    UpdateHandler_6__is_done__q2 <= UpdateHandler_6__is_done__q1;
  end

  assign UpdateHandler_6__is_done__q0 = (UpdateHandler_6__state == 2'b10);

  always @(posedge ap_clk) begin
    UpdateHandler_6__ap_start_global__q1 <= UpdateHandler_6__ap_start_global__q0;
    UpdateHandler_6__ap_start_global__q2 <= UpdateHandler_6__ap_start_global__q1;
  end

  assign UpdateHandler_6__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    UpdateHandler_6__ap_done_global__q1 <= UpdateHandler_6__ap_done_global__q0;
    UpdateHandler_6__ap_done_global__q2 <= UpdateHandler_6__ap_done_global__q1;
  end

  assign UpdateHandler_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~UpdateHandler_6__ap_rst_n__q2) begin
      UpdateHandler_6__state <= 2'b00;
    end else begin
      if(UpdateHandler_6__state == 2'b00) begin
        if(UpdateHandler_6__ap_start_global__q2) begin
          UpdateHandler_6__state <= 2'b01;
        end 
      end 
      if(UpdateHandler_6__state == 2'b01) begin
        if(UpdateHandler_6__ap_ready) begin
          if(UpdateHandler_6__ap_done) begin
            UpdateHandler_6__state <= 2'b10;
          end else begin
            UpdateHandler_6__state <= 2'b11;
          end
        end 
      end 
      if(UpdateHandler_6__state == 2'b11) begin
        if(UpdateHandler_6__ap_done) begin
          UpdateHandler_6__state <= 2'b10;
        end 
      end 
      if(UpdateHandler_6__state == 2'b10) begin
        if(UpdateHandler_6__ap_done_global__q2) begin
          UpdateHandler_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign UpdateHandler_6__ap_start = (UpdateHandler_6__state == 2'b01);

  always @(posedge ap_clk) begin
    UpdateHandler_7___num_partitions__q1 <= UpdateHandler_7___num_partitions__q0;
    UpdateHandler_7___num_partitions__q2 <= UpdateHandler_7___num_partitions__q1;
  end

  assign UpdateHandler_7___num_partitions__q0 = num_partitions;

  always @(posedge ap_clk) begin
    UpdateHandler_7__ap_rst_n__q1 <= UpdateHandler_7__ap_rst_n__q0;
    UpdateHandler_7__ap_rst_n__q2 <= UpdateHandler_7__ap_rst_n__q1;
  end

  assign UpdateHandler_7__ap_rst_n__q0 = ap_rst_n;

  always @(posedge ap_clk) begin
    UpdateHandler_7__is_done__q1 <= UpdateHandler_7__is_done__q0;
    UpdateHandler_7__is_done__q2 <= UpdateHandler_7__is_done__q1;
  end

  assign UpdateHandler_7__is_done__q0 = (UpdateHandler_7__state == 2'b10);

  always @(posedge ap_clk) begin
    UpdateHandler_7__ap_start_global__q1 <= UpdateHandler_7__ap_start_global__q0;
    UpdateHandler_7__ap_start_global__q2 <= UpdateHandler_7__ap_start_global__q1;
  end

  assign UpdateHandler_7__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    UpdateHandler_7__ap_done_global__q1 <= UpdateHandler_7__ap_done_global__q0;
    UpdateHandler_7__ap_done_global__q2 <= UpdateHandler_7__ap_done_global__q1;
  end

  assign UpdateHandler_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~UpdateHandler_7__ap_rst_n__q2) begin
      UpdateHandler_7__state <= 2'b00;
    end else begin
      if(UpdateHandler_7__state == 2'b00) begin
        if(UpdateHandler_7__ap_start_global__q2) begin
          UpdateHandler_7__state <= 2'b01;
        end 
      end 
      if(UpdateHandler_7__state == 2'b01) begin
        if(UpdateHandler_7__ap_ready) begin
          if(UpdateHandler_7__ap_done) begin
            UpdateHandler_7__state <= 2'b10;
          end else begin
            UpdateHandler_7__state <= 2'b11;
          end
        end 
      end 
      if(UpdateHandler_7__state == 2'b11) begin
        if(UpdateHandler_7__ap_done) begin
          UpdateHandler_7__state <= 2'b10;
        end 
      end 
      if(UpdateHandler_7__state == 2'b10) begin
        if(UpdateHandler_7__ap_done_global__q2) begin
          UpdateHandler_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign UpdateHandler_7__ap_start = (UpdateHandler_7__state == 2'b01);

  always @(posedge ap_clk) begin
    updates_0__q1 <= updates_0__q0;
    updates_0__q2 <= updates_0__q1;
  end

  assign updates_0__q0 = updates_0;

  always @(posedge ap_clk) begin
    UpdateMem_0__ap_rst_n__q1 <= UpdateMem_0__ap_rst_n__q0;
    UpdateMem_0__ap_rst_n__q2 <= UpdateMem_0__ap_rst_n__q1;
  end

  assign UpdateMem_0__ap_rst_n__q0 = ap_rst_n;
  assign UpdateMem_0__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    updates_1__q1 <= updates_1__q0;
    updates_1__q2 <= updates_1__q1;
  end

  assign updates_1__q0 = updates_1;

  always @(posedge ap_clk) begin
    UpdateMem_1__ap_rst_n__q1 <= UpdateMem_1__ap_rst_n__q0;
    UpdateMem_1__ap_rst_n__q2 <= UpdateMem_1__ap_rst_n__q1;
  end

  assign UpdateMem_1__ap_rst_n__q0 = ap_rst_n;
  assign UpdateMem_1__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    updates_2__q1 <= updates_2__q0;
    updates_2__q2 <= updates_2__q1;
  end

  assign updates_2__q0 = updates_2;

  always @(posedge ap_clk) begin
    UpdateMem_2__ap_rst_n__q1 <= UpdateMem_2__ap_rst_n__q0;
    UpdateMem_2__ap_rst_n__q2 <= UpdateMem_2__ap_rst_n__q1;
  end

  assign UpdateMem_2__ap_rst_n__q0 = ap_rst_n;
  assign UpdateMem_2__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    updates_3__q1 <= updates_3__q0;
    updates_3__q2 <= updates_3__q1;
  end

  assign updates_3__q0 = updates_3;

  always @(posedge ap_clk) begin
    UpdateMem_3__ap_rst_n__q1 <= UpdateMem_3__ap_rst_n__q0;
    UpdateMem_3__ap_rst_n__q2 <= UpdateMem_3__ap_rst_n__q1;
  end

  assign UpdateMem_3__ap_rst_n__q0 = ap_rst_n;
  assign UpdateMem_3__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    updates_4__q1 <= updates_4__q0;
    updates_4__q2 <= updates_4__q1;
  end

  assign updates_4__q0 = updates_4;

  always @(posedge ap_clk) begin
    UpdateMem_4__ap_rst_n__q1 <= UpdateMem_4__ap_rst_n__q0;
    UpdateMem_4__ap_rst_n__q2 <= UpdateMem_4__ap_rst_n__q1;
  end

  assign UpdateMem_4__ap_rst_n__q0 = ap_rst_n;
  assign UpdateMem_4__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    updates_5__q1 <= updates_5__q0;
    updates_5__q2 <= updates_5__q1;
  end

  assign updates_5__q0 = updates_5;

  always @(posedge ap_clk) begin
    UpdateMem_5__ap_rst_n__q1 <= UpdateMem_5__ap_rst_n__q0;
    UpdateMem_5__ap_rst_n__q2 <= UpdateMem_5__ap_rst_n__q1;
  end

  assign UpdateMem_5__ap_rst_n__q0 = ap_rst_n;
  assign UpdateMem_5__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    updates_6__q1 <= updates_6__q0;
    updates_6__q2 <= updates_6__q1;
  end

  assign updates_6__q0 = updates_6;

  always @(posedge ap_clk) begin
    UpdateMem_6__ap_rst_n__q1 <= UpdateMem_6__ap_rst_n__q0;
    UpdateMem_6__ap_rst_n__q2 <= UpdateMem_6__ap_rst_n__q1;
  end

  assign UpdateMem_6__ap_rst_n__q0 = ap_rst_n;
  assign UpdateMem_6__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    updates_7__q1 <= updates_7__q0;
    updates_7__q2 <= updates_7__q1;
  end

  assign updates_7__q0 = updates_7;

  always @(posedge ap_clk) begin
    UpdateMem_7__ap_rst_n__q1 <= UpdateMem_7__ap_rst_n__q0;
    UpdateMem_7__ap_rst_n__q2 <= UpdateMem_7__ap_rst_n__q1;
  end

  assign UpdateMem_7__ap_rst_n__q0 = ap_rst_n;
  assign UpdateMem_7__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    degrees__q1 <= degrees__q0;
    degrees__q2 <= degrees__q1;
  end

  assign degrees__q0 = degrees;

  always @(posedge ap_clk) begin
    rankings__q1 <= rankings__q0;
    rankings__q2 <= rankings__q1;
  end

  assign rankings__q0 = rankings;

  always @(posedge ap_clk) begin
    tmps__q1 <= tmps__q0;
    tmps__q2 <= tmps__q1;
  end

  assign tmps__q0 = tmps;

  always @(posedge ap_clk) begin
    VertexMem_0__ap_rst_n__q1 <= VertexMem_0__ap_rst_n__q0;
    VertexMem_0__ap_rst_n__q2 <= VertexMem_0__ap_rst_n__q1;
  end

  assign VertexMem_0__ap_rst_n__q0 = ap_rst_n;
  assign VertexMem_0__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    VertexRouterR1_0__ap_rst_n__q1 <= VertexRouterR1_0__ap_rst_n__q0;
    VertexRouterR1_0__ap_rst_n__q2 <= VertexRouterR1_0__ap_rst_n__q1;
  end

  assign VertexRouterR1_0__ap_rst_n__q0 = ap_rst_n;
  assign VertexRouterR1_0__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    VertexRouterR2_0__ap_rst_n__q1 <= VertexRouterR2_0__ap_rst_n__q0;
    VertexRouterR2_0__ap_rst_n__q2 <= VertexRouterR2_0__ap_rst_n__q1;
  end

  assign VertexRouterR2_0__ap_rst_n__q0 = ap_rst_n;
  assign VertexRouterR2_0__ap_start = 1'b1;

  always @(posedge ap_clk) begin
    edges_0__rst__q1 <= edges_0__rst__q0;
    edges_0__rst__q2 <= edges_0__rst__q1;
  end

  assign edges_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    edges_1__rst__q1 <= edges_1__rst__q0;
    edges_1__rst__q2 <= edges_1__rst__q1;
  end

  assign edges_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    edges_2__rst__q1 <= edges_2__rst__q0;
    edges_2__rst__q2 <= edges_2__rst__q1;
  end

  assign edges_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    edges_3__rst__q1 <= edges_3__rst__q0;
    edges_3__rst__q2 <= edges_3__rst__q1;
  end

  assign edges_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    edges_4__rst__q1 <= edges_4__rst__q0;
    edges_4__rst__q2 <= edges_4__rst__q1;
  end

  assign edges_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    edges_5__rst__q1 <= edges_5__rst__q0;
    edges_5__rst__q2 <= edges_5__rst__q1;
  end

  assign edges_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    edges_6__rst__q1 <= edges_6__rst__q0;
    edges_6__rst__q2 <= edges_6__rst__q1;
  end

  assign edges_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    edges_7__rst__q1 <= edges_7__rst__q0;
    edges_7__rst__q2 <= edges_7__rst__q1;
  end

  assign edges_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    updates_0__rst__q1 <= updates_0__rst__q0;
    updates_0__rst__q2 <= updates_0__rst__q1;
  end

  assign updates_0__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    updates_1__rst__q1 <= updates_1__rst__q0;
    updates_1__rst__q2 <= updates_1__rst__q1;
  end

  assign updates_1__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    updates_2__rst__q1 <= updates_2__rst__q0;
    updates_2__rst__q2 <= updates_2__rst__q1;
  end

  assign updates_2__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    updates_3__rst__q1 <= updates_3__rst__q0;
    updates_3__rst__q2 <= updates_3__rst__q1;
  end

  assign updates_3__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    updates_4__rst__q1 <= updates_4__rst__q0;
    updates_4__rst__q2 <= updates_4__rst__q1;
  end

  assign updates_4__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    updates_5__rst__q1 <= updates_5__rst__q0;
    updates_5__rst__q2 <= updates_5__rst__q1;
  end

  assign updates_5__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    updates_6__rst__q1 <= updates_6__rst__q0;
    updates_6__rst__q2 <= updates_6__rst__q1;
  end

  assign updates_6__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    updates_7__rst__q1 <= updates_7__rst__q0;
    updates_7__rst__q2 <= updates_7__rst__q1;
  end

  assign updates_7__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    degrees__rst__q1 <= degrees__rst__q0;
    degrees__rst__q2 <= degrees__rst__q1;
  end

  assign degrees__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    rankings__rst__q1 <= rankings__rst__q0;
    rankings__rst__q2 <= rankings__rst__q1;
  end

  assign rankings__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    tmps__rst__q1 <= tmps__rst__q0;
    tmps__rst__q2 <= tmps__rst__q1;
  end

  assign tmps__rst__q0 = (~ap_rst_n);

  always @(posedge ap_clk) begin
    if(ap_rst_n_inv) begin
      tlp_state <= 2'b00;
    end else begin
      begin
        if(tlp_state == 2'b00) begin
          if(ap_start__q2) begin
            tlp_state <= 2'b01;
          end 
        end 
        if(tlp_state == 2'b01) begin
          if(Control_0__is_done__q2 && ProcElem_0__is_done__q2 && ProcElem_1__is_done__q2 && ProcElem_2__is_done__q2 && ProcElem_3__is_done__q2 && ProcElem_4__is_done__q2 && ProcElem_5__is_done__q2 && ProcElem_6__is_done__q2 && ProcElem_7__is_done__q2 && UpdateHandler_0__is_done__q2 && UpdateHandler_1__is_done__q2 && UpdateHandler_2__is_done__q2 && UpdateHandler_3__is_done__q2 && UpdateHandler_4__is_done__q2 && UpdateHandler_5__is_done__q2 && UpdateHandler_6__is_done__q2 && UpdateHandler_7__is_done__q2) begin
            tlp_state <= 2'b10;
          end 
        end 
        if(tlp_state == 2'b10) begin
          begin
            tlp_state <= 2'b11;
            countdown <= 1'd1;
          end
        end 
        if(tlp_state == 2'b11) begin
          if(countdown == 1'd0) begin
            tlp_state <= 2'b00;
          end else begin
            countdown <= (countdown - 1'd1);
          end
        end 
      end
    end
  end

  assign ap_idle = (tlp_state == 2'b00);
  assign ap_done = ap_done__q2;
  assign ap_ready = ap_done__q0;

  always @(posedge ap_clk) begin
    ap_start__q1 <= ap_start__q0;
    ap_start__q2 <= ap_start__q1;
  end

  assign ap_start__q0 = ap_start;

  always @(posedge ap_clk) begin
    ap_done__q1 <= ap_done__q0;
    ap_done__q2 <= ap_done__q1;
  end

  assign ap_done__q0 = (tlp_state == 2'b10);

endmodule

